PK   c]W����,  f�     cirkitFile.json�][s�8�+[�q!	!�c�jf�k{k�!I��j;�qgf���G������8��<t'��p�>}���A�ӛ�j[��7]��&�br��u�=͂�j�h������.��n���t���?l7z�,R�#%T��X��a��I(t���s�L�"
��]���R�X$a�E/W�p�%EX�
���
�9	f��l)�T�e�G��H�0]*ʒ�"�d$����uvY͌Ո��]�Ǹ��=�uW��)�{�A+[*��2�T��"\F�y*4���L3��E8���Y&0C�����W����ؐ�]�,�B!Y���%̬������!�C��z�4�j�}��$�5H�����l�9�O����Hj�H�č�.II\a.=F�5Fҍ��!���-6а{�!h�Q�,�q�/ ]6G\6*��@ �@.r����{֠q�Ծu��>��:�3ϙ�f#e�^$�Xa�?� u�S0ȿF� �������8�@]5j��oi�̩��3- k]�S������
�T�N}��L�.���a�%�0���ւ/����8rm=���W���F�⃿����DVK���I�-1�I�%!ѢH��$Z�ue�p��H�a4�e4�e4�e4 f4f4f4f�~X5�(X����4-K�s�#���(s��e�i�*�4(4\,ZI�R��P��X���p��A��A��bh��@#th��tT-坶ZY;=.���Q.���NS9��uzEBY�].�&u�ǡ�%��M��8h��4�B8�#h-��LC�*�gZ!9=��b�����gZ�x���r®��-'l����5�����I�-1�I�%!ѢH��$Z2�������������ÌČŜŜ��iP�iP�iP�iP�iP�iP�iP�iP,hP,hP,�B	�Q��	x-���Nj��ZF�\N�k]�r^����	x-��\N�k]��r��:��ZFg\N�k�ip9�et���g-O3����لEU�\�t<V��-��J�j��օ���k��r���?q	~B�|S��G̣���sj���9��lx :�U{�����ԘM��g���p!,b\�̸��S�K�L��a �p|�2`���j�1�U{<�;�-ߩ�[�0;$Q�K��s�����Y���;�02&�� ��߈�
	�Q�/�-��d���iX���L�o
WJvml����֞�g�{�gx�Y�I�ee���]Vɳ��?.�#dF�Z���q�4 �.NY �>�Gv�7 �d�W2��� �M��;���a�J@{�`1�6 Y����Hn[|"� Y��[�E��2rF1����)�1@��.g�Z5���C��rH�֮.G����(Z�"�U����2���gN��U�?N�qY��z�u��6/^��>oQ���U���uP٦Q�@n����1��D�O��������/K��ð�dXD�{z+����Pa1ʰ eX���zc�z����'��og��C�&���ӜcAͱ<�nj�]��ȱ��XP�;zW�	8���M(_�%_ိ'C��h@��bLC`�X`a+��'��y����`����ӆ}M�:��؃�6`��C�����9�+x�CO�=
=m�[���B��a*��cJ=�p�K�v	P��&`@o�����P�f�����U�g�e_<i'�2�9k��d;ǖ_,-|,u��ά$��m�Yaf������3ۡ-�US��=��������m����mn{ۣ-y��ۣ�'&la{����ս8�	B��1!�v�ct0y|�G����&y�;ǋ��{������J!���%���{fu�K�w�b�)��!��ޓ�q���Z�܎{�0&"�=<tɸ�TcI�S�à�}�~��Ž���(c@ԇ������g���I�aƋ� �F�k4����|��6(��������Y�5EǦh�ďM|�$�Mb���a�<6�aSrlJ�M�ؤ�M�)6eǦl�Ğ/��b�/_��Z��r�����r�XW���j�U��r�4�f�Y$�.�(_�I�3Vf|��Y\����/�b�˦��*o�뻿�Mn�}o}���n*m#w����jگ�^�,�se�<^��1ͻ�n4[�P��[ťY�eJaL^	�rU$aQ��X�E��9���|�:��
�`[W���`YPl7�પWk}��k�dʢ�𣒙����Tv���uTJ��x�9�g�#Ż�S;�Xͱ���3|R)�r,�
J�=��������2ճ�����e=u�!9șQ
r�F�(cص��q���P��});���ņ�v��C�:��w^��N�>�gL\�wA�9q�^{���>�}����^p�A��W�|�`��k�;o[���j�6������Q��ٜ�8�W�T��~:&��/C%;�'l	Pqf"�8OåXf��)�:���u���-}w�8#����1n�������; �s������#��`��\=�?�f��C͞),QءU� C-����8V�t��M��+��J"o�����=M�LPp����ٱ7����6?�A����o�:�����ߟ?�f���7�	���n��y�7�9�*��N�Ɲ��v�r�_������f�f`��}���}��S&�{���C^�������^�*JY���Y9�n����H��5�n�L�e��,59�ȵy�D*��lo]��
����̢�:�¬�����U���'��E?���ό�t��p����3��j���2���`*��0�M�S1/eYh��>n@�n���9��� ��¤�Ex���X�)�v�)Z5[3ށ�$�<�Y{���CͱX�y"������*X&�9���;]�|gEc��������u��{N��N�^��/�n��~����vr�>�	�~�W7��?�	f7by�|�6?m���)ZezS�T�mѪ��ǯ��}����a[m�/ys���~ssت���m��.۝=zum�=��a�d`%f1���[�g����M�d� Ǆ1���6��)�M���L�]�#&�S����<�h�� f��9:p�I���
�,�h����d�9�=)��\R��(�ٱ�&u�^"�M�1���D�!6�c�`�D���Ӵag�ݢ Pj�8<k�C�b1!�)b�iYL��b��D�R&�v;�� ���Yv��@)0�M�ٔ�'a����)��gERc5e�a ��[�J����N�f	�Q�d	)���%cNg��T�_���8C���|��O�s%�Bo<=D�=LA�	$�Ä�i��������!g�(�E�^T
ȩ��$,�dĤ*i� �Y�A�ܞg H���Q�$hL0��,��5�4��`�޽u��F�=TJ��t�!&�.&�F���E{7{�5zR<�dy���b��1����Y��$�M� ��,$���	�M�-�fjڼQ¤�E�<�_'-c��e���ep�l�y��!ٮ�?�)
)��z�9�b�O]S:N�{�b�&�F�8ς�� �ٻ1��I*�rL�Cx
Ğ�,�9	fS���&��&▄��{�al������ �I���{�KARp���`�	��Ex{����(�b�T6�A7ɻR"rJ�~@B�R�C��!`��S�2M�md���2��3\n���] � K�&���c&|�m<����|��Y7|���3|ʲT�|AX��T��F����ك'>���(�r�r�^.�]W�z\Y��?�����|��ן��?4�~gM�}
�~PK   c]W ��!�} $� /   images/c261b03e-8211-44a8-b3b9-e5822ea41eae.pngTzPM�6��n�����ŃY,��I�`��;dqXdq<w��~���޿����g�F�9�tw���26����.b�߶���w��«��		(�!ט��d�� /��*/O�����d��%苤ʠ6Q��i�.;�7��w��$�5 V�Hm��#ˋi���%"uȨ!$�8ܰ.���Mܘ��Ԣ�4_]{���G�Ӽ��[���J;-m���%)rܽ�H�� �T�kQ�w�Ak�#���&/zn��1����!������oj8ن��QU��{-�
Ø��%��?�_�[�$mn*$�-�����o��o6�m�?En��5�{U�4�0���'aT5��3�K�y��IQg6DN�¬���u���y�ؾJ�!�D��i{�CA��d0�֛���)�G�N��e�Jj.$,"�"��:"�Oh!���������	=l�X���>.'�Rp�ـ$�zZ���?=:��%{i�_?�
͐��������?GAwy��t7c88L�<\v.��ATOUE�}j�����pptp�
���+��WS���nq�GK��C�PPe�[���b�1��S��zc*�6.�����~���Ҏx�;�lb2%R�cE��C��ݯ��9:���ʄ�p荳XM��}�}�,>���+��m�lb����G��E������X�w����3]D�� !Ƅ�^;e�!G�d$; S4d��q:��H~��Tik�+^t;�[<����:�;<�w����-����'�ӦzL�|�G�O�OcW9�T�I���6��������|�����~ZV^��N�Z�&�([؊��Pkj�,`BI`û�	ŉK�Ѩ�O�n�6G�jTuT�}F׭�#�7�MA:���ڰ q��ej���V�j�?�+�r=�z�_^�A� M�u��o���@����W���N�2L2��v�����	���\^���T
�D����:��;X���g��P��Y1 �w�� ��2�Z||$Rsd��[��xx�r��xrht�e(?���r���Y^�T�#l�o�h_���%��r
�4���!6Θ�$�r�\X��p�V�l���T
k:f�������e�/�V_,��J�t��;ϼ]-�I\�+ζ�?�i�����|��=?Z��ẖ�K72İ+�-Emq��T�d�� ��wt�����<R���LEC�JJܬ(k,bҗ�Q�2a�L���0��(Z�@Ʌ����9�e?MS�
�#b�q�J�0��Z�������`�}5���ZQ�&P�~{p��	�X &Z��'dn��j#7ժF����Pٜ�i�e��5��9��tf����@��Cz��׎Xx0t�j��B�w���(?����&N��1p�2r���ǹ��\�'/=����zM�uuMg��?D���!DXE��
S��^�9��~�'*}��S&LJN&Od����K���<8C����\&���Μh�1�q�(���3�m�8V�����X9�ā�D���[���E�xz$ȭs|%��M�j�-r� ����B���KRJ��lOɑ���#r�N�5���`�C+(,b%�ܑ���p>-���?G��R�=�]^^��|�K���6��}�	�����_�eM��:m�M8נ���=��we,�O�~��Oz<��ZIJw��u���:� ;��F����+�����'tp��x�ۙ�
!K�-c�l������#�Ӻi�qӍ�	�F4����:1H���#yXц��M���p:F��`���* l�J�`����ɻ�8<r�0S��!R2^5z/�[�{��3�ɪ�(I�l%ZF]���[r�Nu���F�Cj�&�~G���Φ��R"��*�T�:td����F�h xv��MC�[��)�P�F�J5�NK'�<�L��u3`��f'0+��d_D+��������(�!��H5�1��x��κk�L6��V�'�%�/�![���*5����6`���1��I��������<y��^��Ϡ�6�h��&5T�IL ���A	��N�D�m�/�)G�f���x�V�,��ێ�h�� �U`6G��0";k��F�~���|��Q����v76�T@PsHKj����!����Ӆ�u�͍	]Wrt���Yf�"�+W�~�ƍ��6v�Fj��($߅X�)�ˠ�o�u,!r�r��kTE�,������3��kx^]�'$8����Ifw(~�.���_������i�p��si��b�{�������h<�O~�Ġ��}�k��*���$X�ۏG��ߧ��ض�?�~��1�����y;!�63�X�u[�����LqJg�1��N�p��Ui����G'�j���}�����̕ ��%�\z�}�<Yj���$I�11<�ܼ*:� kq&K:�^��]����"�f,����rO��ڛ�ve4�DY�ĺG2s�^�q�Q�V���_z�ckdF�1�9�9q�����ot�V+{]��R0S.jvT�5ꇠ�޻ZKgYk.����6�I�!l�H
q�?5��ж���q=!C[I��M\�弈�x]������۷|/Z<�vʁa�% ~m�Ƅ}�ܖ�M�s�d�Dy��`�@�]�X�I]ZG\h:�S̜f�
�����
Qi>uZp+7Yu@
��s�4��?!i���i��17� ZZRK#g�!-��E�/�ni��K-��
�����0.h��5��R�_�ֿCi��'���*D�K�3*(�f�m@SB�'.�9�G8Oz�A`����Qm���|]t� ru�8>"�v=9�5��^��U[������z�@X��n�<�{+)�������6��Nz
���(mR�BLV�t6+!�-�Ne�<�3�B��'���A�ۮHNҎP�(4c��)�s]��Vn"ʘT<�'+���6
v�m�"2CVͤ%o�s=�hZ�8b��Չx�~�V��{J#����a�Jjø��PL�o��C�[O��п��1L�M�D�qX_�α
`piwb��s��"q�GM�F��X����j0͢" ��w���0'�h*�\@�lkZ��i�>����nj��z��ڀ� ]R��/�o�j��E�?�#<���_X�	#\t��w�b�ڵ����X';o-���l�ɸ��9g/��lT�#=�K��X��Z�3Z6�N���w2��j��XEN�ډ��s2E��Yt�$�m+e�}���Ɖ�x:\%�ZfR�sj�_�{��@+r�ы T�(���M�~7���y�Y�4[r�Y�ں1oM}=�bE� ?~�������!\�;�E���Z;��q%RpJ���P��E�)�E��AT��R0{X�ȠJ�-II�p�1�/s��IH���}j�k.��1��%�$���8-ֻyPB1�{�,��;.�q���j�?@��t6V�{E�nAK�����ǣ~OՔ��Mԡ��j �k)˄���u���4Rb��#`^6KH-���PbR4G�+�t�C��1��nK�i(��j
Q-�@�$	�:�C8�5a�[9m�����b��$6X�bm�Myx�r����Ia5Y��N�1�U�¼�xn�
�y�"�Ɣ
&;�"R��>�Y���uOA���ז���B����ݠ�[�Z��a��}ݻ�Dka��?['uH-^�kFk�|�f{y#u�)Xd�(.{4IsT�(W�;��8�:��䅧RU��\�!��ʊ>�l�Ģ���($��|t+����rM��X
f��������p���"=e�W��[v.�C��٤�;d��_~�J6a!X?�xЈ~��!g�}�g;���uҾ��5����.e��Z�Kk�S��Q��n�]�u9|���[j�.�h����w�&z=<���pR�U�����5��Cv��Q$U�ËX9gRe>�Vӻ�'�|¤E���\���Z���+�S��;�̧�<$s�;� ¶�w5� �od[�\�П]��9U^�1�J���hcQ����{����>w���L�>�f���og�	8tC�$���)$���MLܒ�W��P�d�gWL��	X�zBQ������j��Gx�r��ʪ��ݜ)u]���ٜ�A{Oۤ~G�u�ݣ �b�����^_������A�~�n�Ã��f����p�����v\`�X�,�6 �p�-�I������ϵ��J[�#��Ԝ�T�n�t����&��7y}tɷ���͢Nm�#�k�����~G� ��s�@��B�-b�z��m[6��i�R�>Ĥ]��9L1��x%W�Z�r��pb5t�%o�Qek
2�脃N����'6���@�����}O�"��ƙ�7b냲Ϳ>C�,���(>!W`���܈�q����Q*N����<� R*J�	-��X��75�)�����g��_ĵ��
h�JK�G���4�ڒ��[�$S/,.~o��6)9B���!���P��Ǵ�?��U��7}-�� �ݛ~�)���S���E���O�%�D�?�~�E���\
����s 0C�����JėF"v%a�����"��lv��]x���:��:���?܊:s����DF
�D���V�6�,���~�s#��w�m����Q;7������� �Kw��~m��h�l�H��ِU�](fk����]�۱ܡ��h��5C3cS�0�l�18ָ���H�įB�c��P��V��c�8PB)�&�;�a�J�ܺ���U{talΙIw�'̻���i�O�ؕ��˞��G��YB%��EaUܰ�Z�$���j�ԭ�"Q�ԫD�Vif>����ڥ�"a���x�����	-\����5א�� ��^pf����]L���,�=	)�-Fn�� v�@2�D+��My�; PC�ۦ�--�?L+��1�,M��k0>V�-d�QH��G�<mR�*뤈v�-��vb�x�,G�-k7eV�<�Tg?�z�ct�
S�0r :��<Zu���8��
��/p���*��W8Z&��|�R%`\�Xb�bJJ��/R�}���� �~��\v��ܸ���=h��B���hq-���sc�Ɠ�-vA>�9�.���{�� '('��l�5��vQ}�i�OIT&l("c� �`���ZME�T��q�'*����)3e��3S|��/L�3���Ư�?�����t:��C�^��|�2{�v�-.���N��ڥ�^X5����<d�����_a���1a�74�4bb�n��E�/�t�WE� !�!:a�`���@���b��aՔ��ŨAe^3��)��ZD�/���M�lcM��(���ȃSa�Ru������p�`�}t���]pS�T���(ǹ0��[����N�����:muĨ�|��w���Ua�(�s��;�1�6�#L1�·2���蔔(gajj�A�H>�g����_�"t����C-Q�������4_�zһ =y��J//�t�ZC/{����>1S�;ʷ|��_�=.�#��,��3�	8ϛ�[�<�}�<�C{&&P�H�`f�~�����,j⿬{P�jx�{�.1���S�h���0KTꏈ�bB؈���W�L���O�"r>�/D�ϟ��Q��Zc���I��̚��-<e��&����J��'����a[��=I�'O[����� @+q3�,�[������=�J(_�ߦ���Z@�~���AIO,��Z6�� �jwU���T*�����*��=X����9c+=���X�nAou�zLm$����>�}/�
a���w�{�qgj�.}����3ehP��Uyk�h*Ko���^��'8��i�"E�����8�z<�a�n����:��2�2�R�����u*��GRD�n6%��7Mr���߮��h@K5J��/�PA�Ab��v�uJ��Pj�x��w������q��ˀ���g����q���*��o���B5aq��]��J���G'��jb?����$_���J�w��5K�E�A�0�ܬ8�)pF13J4���u'F�3��4!WP^�a@
�Ai�v�k�B�_C6�7�
�3c*���udU.�ՠ�f��G2|�����A4��[Ʉu����&���X2����^/�R�����ŖNl��@�k�B���DV�I��m9K��l�A�_U5��3j�3��I�_��7�}�#� s9J�h��y��{�wBP�A��ȥ�P3�X����o�m�}�Dl�ѻT҃�ȴ�58����t�3��岿����:��� t�P�nz/�����ep�T�7���C�@�R6��{��р{Ez����Z�@��h�ZЯq��h����i�)�� �Y�@���-7NH�;�ޝ,�������mW�]�����Z bpEg��5�]'�����������R��i)~x\�z?��7�|�Tei�Cn_P!�[���+6m���8Z����}A��y����"7����Kb��ô@'��p����l�-�j)���@B�PzjIE�kG��F�0C1�A!SӸ27���K��\��=?�b e�g�	��i=��<h;lD�j���b��q~�ͼ�Z�w��j;�z(���NB�fgH:���O~�x0L������D�ź��B6�ե�®�!�-���I�*��l��e7M%��ȫ��*o	����p9���#n�t�㈃��ɰ���Q��v���d�r�&��gX]\�dY�&��`��2�� �1�p�Je�Qj�#^��P`��$.\c�(:��4��xɈ�}.|��,���ӁR4��6����l���;G���'�s���>	��#�`p�4�m)n5�й�V��a7��㣇�Y��%���w���rR�n`��gڟ����Y�n�יĝ�`Lζ�Q�R]\�5��I��ݒ��c���&�X�HY�"i��-�vPD��Vf(j�5Tf��߈���v���nG��:`����4]#�US��?
��	���q�1l;Us� }TkkLbW�����0~9��KV��'�{��V<��0(�7�׫`�b�D!�F�f�� �a��ۻ�8�<�]@�v�t�\�����
(Lg��!js�{�h�Q��@�D��d-6�>�����zQ�
okT����	M�+�M���+!���_X���(d��d?f��H��'a�����ע�	������u���7��ʎ�r0%Q�y�c�ĎWis%o�Z�+D��U6�f��$h�s�3�Y�į?,�
���Y�d�M??�mO?��+��.�|1�İgh���S*-��rt�|�
�o���
U�Z$�/��Ȏm<��x�|Y�}��9�s��3$��Q�вg/ْi�gwY�;z�x䕛
6$(\��//Fʱ)0�E`�9���c@QM�:����3�2ȃdew��`\�D����<s䟆�Pk��dU����qZi��Oô�z�DBDr1A\��7���Ub�2[q��>�䏧k�Z{��. E��C�_0�>o���^?B���Ae,TyPFXݪ��Z~��Ƃ�a�����H�X~�o���z��m)�\d6*	���BS��5�T�R�r�ho�'o����G7ވ(f=��> ��r}e_8�Jz՘Ũfh���«osV�O.�V�������-��k�o���H��ٻ��c��c*�l*~a���c��`)�F��9��#QL�z��R���N�L!�M�Wx��ՌĤ]����haô��m�Wq�^����O�Cv����O����Y����5����ϭK����-����~gK3�;�`K��OE��?�I��}4wH���	Z�rw����!��v������d��8��o>�E;���*�����99�H�/���e�FX�Zsw y}��}�f��(�����j�s�R�;��i����2�d�;�W@a�G��g#��0f0��n�[�I�OVN�R���1h�w�V�L�M�[30Uk1����m��ܥ�ܸ��jY0�ܼ���	Qi�B�*2=�q��OVxX8�Ƚ+ ��@���/WɯY�BL���'�[{'@c����P�I��)J,P\�vӊ���beUhs3?5���WF]I��ѿ���Q��_k�gx���uL,/�uO��H�ؿ��gk��$~ņ�ۼ>�Mi�s�b�{��h\�b�g�����R�e�~Y<$�ɓƜj���s�<�켒����^b-�bZ���3�oa��������ec�Iӭ��_%^�Bz��,6���us�J�#u���ϓ���\e��!z��?n�wq�e�F�e���"����0r�<
�p��'��o��'@=���r�B�R��r�u<kS�V���C		�͕5�_짬�UmUU|�^�F�:,j�Qu�ud�:^���M�CM$��:�PV�]�!�^�����`W&t����x.�3��xw �'�>����аg�����F�D��ɋ��X,�~��?/[���/	��|���y~	�\þ�e8-����ֈK���߽ p,��#�]Q�H>�7fY:�(���G `��/�C{�)���:�q��W5��Q�'4w���S���/���(s��V�5{w��*�CT�5�-�����l<��{��zz���O��.$�3�~�\����"@l&�ۦ붯�>??Gs�xD
z�o�i�0�jj�_�_�r�$����H�r>s���i&���%�Xt���V����':&�n�����&(�I#����x�+T�)H����.�E]|���k�_��vrr�AK��F����L���� ���H1���X��f=�D񐉢#�w�i-�
Y��U����z��gC�f��fR2y�ȸ]3"�Q"��8H�P�j����R	lək]<���) ��[��t����[�)_��DfU�m����Mv�n��V���P>���}���T0/M����ē�f���ͭbB��M���p�F}V�x�T�{���1_���l�G�'0yS�@?ΒPNR��ގ��.��ah�����Y�/�V( 0�͌�9��~6Q���0"`��ߌK���#���!0)����dS�S����і�|�	y�xY�<t�/�"��u�("�~�-���6~�$��>�cN��t�^B9ߓ������t�A�_<�N{�����uk�q������s�55�	$�!�7�0�(ˬ������!��;@e��B�A��[��5t�F��K�s�i��D��u%������
�ZS���7xq���1L��y�Sv�6f��$ĦK�K��MR03��ط��52�uL��.�[q�������Ջ���H�/�������s��M�,v���6Aga�N��w�ӘA�TJ]J��l^]E�������t�=yLz���MO���!Oc�7s|}���7YC�%����o��������j̲J���7�P.�k�So^=�����P-jv��������,z$��I���NP��Y9X�`�k.�DP�p��j�ͨ�+B' ���e#�_�1RBY�p��l��-�n�^�`�,�6l�㢈NU�_5��mp���]c�Sq�&$����@������־��T��8���пb���;fU�*�E�����<a7YT���u��$L4'Y� *&j'����������-0����� ��� �cUikuy��\��LPN�<���4c1�Vjb�z�0:�GZb�$�2���V_RZyz#�Y�X��T:�s����ǫ"�z3�5��W�U[�q�w`/G�J�P=_����E��k���,�������阍��j�lK"�����s�	05w����S�F���e8'B�4�ͷT����ߴl\��t� �*Q�Z���b�*~M��c���)1�b�ɭ}[B9�
�B*=�wJg��'*�����!� ��vT�[��B���.���w;cj�W�s�RC.l��H2��˥3�w6~{x��;+J`�)�H���2�G���(��sn+{v> ֑r�;>�e���Ɓ4R�h&|4~�n}ʴA
:��\c)�?�~?ո�I��r�o���ő�"3:�|z��&�E}�����c�l�..�X�9������yV��_`V:�{�NB�g�`T� ��R^�%�)���t��p�rqꔂ�?3�.�R�S�n��m=��.�q�"����Z�P�|!�6P?E�]&r'�@�P��j�\������٘����e�N6l�/���F����8����ʡ\�k?�V#�~�50�!�����~}�����~y|4�ǇQ	#N�����nܯ�ȴ���N�]��&�珠]%��D�Bxӊ�A7'��R|�/B��9E �i|�5C��8��h��Y5�b�ķ�)dB�H����c7��'�zuSJ3dyv�_���n��~Aӹ�n�7g�z���/�/ۗ����夷(�u��w���7��  9Is#�; �5:z~�'����ް��p����(M�h�;Q�ٳte��z�&����@�rB��d垣TZ�a��1h�S~��M�ɏ�z���I�CN&#M�b|�N�[n��ag���w-�,�B���k�r.8�Lm�;Ɯ���{�3�D���.����_P7����1�{A� �������iT��+E˗3���1bH��XP�|UL;,�K|�z���C4����j���_ڮ�q��MxI���7������T@�Z�6ʩ��в�����"��O'	3���+I��×
��"�9o��>�k�:�X���K�P�ը�� Q5�Z�!"���C5���ƷK�66.s?�As|,�Z�UJ2l�I�6�����r0+��A��.E&��Y{��|{"ĉ�u�ݰY��������PR�+U�w�_Ճ�͍�E��� ��h��̪���2�2ѝL��+e- ������i��H&\o6P���Yn�x��z�d�t��^��\f�#I��Z�p%�>]i�k��ǽxuU����`}��b��5)�����=a�u��#��m������g�ʬ��pW�������9}��*}������}co2�Ɇ*�v̰��'�"��`��;��x+J�(J��E��jʢ��E��ǎ����4)Ԩ�`��8 V�(n�^�h��+.=����͙�QBz��!~+i�gL]:�,e/�F
L`'���<|.
#�j�y�ǰ �d�͌evx9��$�
�]�l���n-X�YX�Ok�����_	�{A�����j�Ǉ�`�R#��|Q�ٟ��k��L��`�#�q���]���A�jM
�M��H`c_��XBT���̈́�D���z�s��f�Iw����7�+.�������G�L3��o�Dw��?>��'�U&�Uq�G�b���{α��ӲVs�}p�=��1�K��9?Ă[�3g:�q"���/��܄��~*�@4NQ��/f����*�}m�I�tM�Ӿ�s�ʹv$��B�n�c|}�F����x2}z��D�AJP��"ʲ�=�F��^^^y�E��&E�gB��3[m�:��(�P�TN���ݸ"�~jjs�/��*	�x�r����K�-��
���"?*"3���*&Ye�-�^�\N����}��s�+� ���k�]/�5��Xʼ�~���t���|����j�㎘~-">_&�ؘ��L���|	�K�3�o0[��L#��$��~ �[��D��@�0@*؊�+�L�t)kz�g1������h�w``��t�ӘV��)���CBp�ҟ�D���5�a�ǾC�����7���E,���Tf�JS� ����{�ӞK���L���d�?�9�XID�� r��p��F�6\�s3�X���_���D�� _w�⚪X�RF���4Vre��VLr}8I�j�$by���@hm㣑�����!5�,8Xi3.�hJ�����E�<@��L�u�3��GpC�O�<XŰ{֐���$���'��zb��TÔغᵽ�Z
�y�����U�]���xۈ�B�o��I�����|�s��R8Y����3�/�yܯG�on�w/Z� w������f�^�}�����׆��?u|�˂�����?'�;xM���ٟ�%����(�3�li@b}��{�+Px�;ř���Q��ݪ�t�"4��Q��$b��f��S�3�C<�J������g%����������/AV'&~��r7���F���Y���<l遨�+����D��:#�q�i��d�� ��J��xIUYи��fzb]� k�V!. _]h���>�9�Z 凍�]
�/�g|���D^]7�e� �;�J�<����4�#.e�j
���
�?�c��}"7>T���\�I� �����,����"�n�%�$���x����n����LQqIy	����e�1�F/��ˤ"��*��R��!��F���Q'�,���/�*�����.[9v��R���!���DG�o��o�[Zq�iWQ�8ќW�/$=��L�<`�j�����q�4�E�D,[�J���s/��Ϗd�N�1�A����Z�OG�zX�H��#-#�}����@�'B9{Y��v�qQ�oUU�+�g�:0  �s��5��Iks�4�6�֣�mؙDݠ����`Z��K�����@~ȹb�:D1�&|-o��X57`E�����[9�5W�,�t��Ǐ��f�����+�Y��6ӫEƹ�K�e��ck�݉%V�A��9bE�u�P����;ޙK=d����X�&=��qa�����v;zu8���ٓ�Ù�A�<A�c����A�,'��r�塀�7:Z������}y��}�ǥ�PXN#��}[��/�4K��#~�}��t}�&�I��A|,n��N/�j�$�s��LӍ������xr�}F����]n<���&!��u)eŔP"W�Bx�;L��]m�Q�!P�?v���iu���������n����y��xug~2�Ӑ��<�_6.��DP������"�?���g�+�5�����w�^�:��~�ȋ�̹?eO�TH�D3_�Hϰ�u��$d����)�v�jDx3&��N�Q��T�(;q�:e�ûp}��暆�}���8�B�����MΗ�6�%���Pr��o:q�c&F�c)� ��	���������V�m
 ��.�1aE����qn��P��ư��ʮ�0��d�av?�X�{��S�y޹��p�I����I�?���[c��J���$o+V�Hc"�l��ΰ��C�lu�}�
�{� �������A6�����u"��{%O�Yp�d�a­4d�W`wBx��k��ZI��Wu�#?j����G-=�W�S�ކi��z�8��$Νd^2ku�Vy�����u�x���P#�,�I(Uꃆo�� *�Tq!�fÖB�<{�>C��6�s����;��]i[ vM�5'K�S�ڵ����鳫�7��7
���q�W>�e��uq�?�!�ү�!W$;�D�X��2�W�g�gG�h$67��/����f��}�	wD���FM�p�5���Q��2e�-���02.9�	u�,ؤ��v+ٓ}h���6�K}�A��y��2�(�
�%YE��ji<�!p�m�xT����!���M>�`�C��=�l��$7?��(�J,���>����w}�zF�]�}��5�=���o�{p�.�`TU��/(g�9g�>��迳ȧW���|�B#@0�O�Z���)fjqN�x*X �g�:�e2�l�}P?+��L�`5i$&��~fW�zDL"��%��?���s'qk�n�On�^�,Kow)�^/kİ
uI�W0��'�_��	O<���FmK+��Sy)6�,$�� �z
�����؂N'�'�ǈ��,���P��kA<��?�A����k5��z�{{(�b�V|����ѴR���ʹ��/#������ei2m�J!y[P&��^��j�*�J�ї�k�bv9bJS?�W�b��ܺ���Opˀ��p��S"��i�SY�R1O��>W��0?ݾ���?^��~�L|��g�vA��m�~B��rZv���/��&�p�`m������$�a�!�O�O�/l!��wY��!�Ԇ�ZTZ���_����e�o���[/�(�5L��Ԙ⦦���F�T��č������Y��g	�b�hh�0Y�ߐ���^�r��=!� �ƺ|AR���cq0U���m�����߂ǳx��z����\��[l������L+�<mNG4q�J�����|^Q�;R�������7X�0NU�UJJ�䯉��6J`�*����8���E��L��ԟ%��)�a�����O�
��Rﻥ���z�5-Զ�#JJ�M?D�����+��,о���/�@q��� ����������zy��W�b"|k��%��.E��H�*d����-;�Z3����ع�Es��w��kZ��Y�|�j�_#�U�GXm�Ŝ����~�ŌT$9sW4��(��S��<�}����M7���7~l�۞���O�cm�a����g������2���7���7&�U���qG�j�M yUf�<�����K�U���7�?�Z�u��߲*5�`G �j�F�bJ��D��=��IR� ~\���-69,��ͻ~������?x`������N�gm��I�9�wc�T������m�}�BUN66�����։�;�0�g��(��m]G�_�p�5�#��S��.�����N���6o?���G���zƎOD�_��t����t~��P�KN�Dm���<�2S���������jƊ����G�P8<SxV��6S����@��u9 <�L�I�iA��z��K���܍��]�R�^���)F��SA�X�e}�Zvͱ��5%fw����O��w��r�l�e}$q+7|��Jy�������P(t��{��%S��A;�nnn6����L��{�;6>11��·����\XD���4�TR=�6R�A�]|��Ga��"����8�Y�X��ϧ�?-�B�?�O#&��;"����՗7�8@�V�x�c[-=�NO��L�M�D�8O.�	ǫ(��a֧����4�rX�Q�_f�������L�bLɔ�����ىkWk��|��?�Ȼv:	3����r���D��x��{��z�<`�to�Zc����w^sŪ�>Z�)-�"���] &byy$pƁj���]���V:$�SLC*�M*,��:*:��W���Aa4������A�Ud�Y Q#52i=��q���yN}3d����̋\�������2J�G�JY�N���r��mWĥt5q"�<�ֈi�"T�x�E��[�����5�ecg��}i�0H��H��ß,՗�%=h (�����`a��1�)�h�K;X�[̬?��G�j�B�0�۔�\?W�=�D�s�3,������Ř|S<վ���ӽGص�k�O=�,2q� @G�}�Ĩ����'1�&�����{t����`Мx�ae��R��y|�iל�R��o9�*��J2�|�Ј��X����B�d2��fʛ�Av8v>�Q�aJ�F�c�w��+���eK��*3�N�Og���7Ǎ]8a�.��9���;"			5�;��b'0�i|��(s�<���먣���E�#�ٯK7�3���Cߞ5��ϙc�A��U^>��o^��S��m���k7�_�M�?�H>�����.�^Q%�'W4޲�@6��Q��)N4V�|.q>� c���{k�K]�T�V���
��8.XB|��#$��
�(��,le�k�}\Yy��>s�2Av���1V�ղ�E1O!74m4֢����L��ܮ���U��y&�s�UB��Z�� ̘��Kߵ������=�i�����[�t���1��<R��H�Qz�X��MX����,=I��9�+�M�t��v;6qr�o���YYE`�����@��H�7rj�$�q��T��0r��B,ކ˛��oIg�%��:��]`�o�1����͸�9���oᘤ�-A��S�Y��&݃��ߤ8J)��1��S�
�o~��۔;Pp�r7w@��x/��Z��=2���9Y%<�}�#��rom�A��/; 0���w����s�s�"����R��Q�C��(
A��Y��?Ͽ1���n�����c������`>5!����gq�����V�N�ƾ��q�Ρ�,�j�	G�X�0�n��J89,��t�$&��A3����c-��N��Ɂ�4.�k�q��v�$#���o]�͓�q�����I�A�ܖ�4�pSY"٧OY��O�y{S|�c�t/���p-'�@(Q"��Z��:���S��	ϳ�X�t��m�Gĩ��ˌO���hTڱ�w�?^��(P�
f�9����З)%%��1R�?fT�
VtYd�[g[�?_7�A�����H�
�+Z�v�[��!иww����4�;�܃h��]��^���>�u>̇5k��j�B8�8p�˶ת�*�6��	��jf�N<N��>��U4v⫐ϊ��jcH�.d��*`n�@���d��Yڟ���#���~�<5abz*r*$7B������@bS���ژi��'_ԧ(.t`�Qf�^��/N����H�D�Bp�� L ����D-�R����z��bx��0�"�w�0LX�D{S���5�H3��vM�������;e�8�xw�2>ql]�T�e"OP�M�p�y���"U4�:2^0,s���B厴�����5]KO�p�!i� ��`6�d��f^C��#;��"B�b�_y5Z�[��}�
_O��{�x�F�"����e�<S���G7Gw����X^w�s�P$i�t�F<�w��R8A��zǛ�"��y=\�/��C��R�T^������ۣ�2$?t�� Q�����Ȫjp��:%���\ճD������o?\s�)Q�Ǖ����� '�����F��O�flGH�uo?���ů�jԆ�?��@9�RrVNả�
dʻ�9յӮ��f�\��E�[�D��B�|�v͌u��"����N166@1��n���[�
h��W����بM���=Ӥ����ܰB�g�St�c�\w���l��E�E��Vb�\[5�ZhyZ����Y��Ƨn�q��S�@� @E�_�������>O���9
�����Áf�Xd�4�KA��j�@Բ7���`[󪡵88ٯ3�}܏PY�q&��R�:����ن�E���� i�%������ʖxxD,��<:�6=����v��&\�:����p7��TJ`XO�wݞ,<+'��8&2�$��wbˀ��q�F7�~l��DKb0t��Y�k�YR���-����=I�I�'X Π0�04�W�Qr�NP��p_>�#��OZ��@��R�%˔_�al�/�.���O�ٷD!�ތ�-���F5%�]n�@�~�3@Bml�߲Á��.����?��T7�_:'ZNV��7�9\g<,���v�.�a֪��a��FD�`�ɪF���P��U|��������Fz=�/��viX��Xa��ժ�ux��7�~V���T<�E�#���~���,����Ͼ�����PUN5�yԚ\�՟���쟁�*��+I0؈��*

�� �t���G��Ôd<��F�,��A�䘼W[�9Z>$st�|8C,���~�m �����k�j�@�hz���sFV/{�=�ͭ�?��K5S���s#��&���2y�'�*�SK�P�����{D=�d�H����B�~&�nI�x`�m$�����9�,��NX���FVk�e�f �����%E̩�*����g�>����6.ߤ��*��N��g|#0���u��Z��ئlzO�Qr�<�_�h6}	kfK�����V<�NN(�����BHᝫ�0���V�-*e0`�'Jl�[������R4���.U�Ú��03���F�Kj���5�Z<��ʺ��T��w.������O=IC�ބ(�����[s�T�
�5��n_s�I�`�~t��E|d�g�n�~s���6��+R]�˞@��F -��g�uI����D,gF���*��ԝ=g�����u�-��Q�F����P$:�Ae���iF��f0����|O�!W����uˋ�lx ��ك�[��°��$�:y�	�&�&w|W�
Q�LfL��z������b�Q�]M�syYf/˸TŪĲ0��/�?��������|"`���iC�:���w.x	�<0��6��i_Y��*�G����1h�Y<O�ٕ�W(Պ��5J���w��>|ۙEM=��@�8m����]N¦�S��լ��12��hr�s�zq1A=벐���k������m�~�rjDZ��������D&z�F�t�%���Τ
D�"�b(v��������,�Q�v=*Y��%�?�%�vż���=[P?�RF.��"��5'{�!h�:��!�uy�ynx������Ą#)<g��{Xߝ��0�s��Jt6��a�G�	!#�9��JY��I,�I��1ͅ(, 

�A�I)wh*?Y�\�-nB��U
�k��� \�bP�*y�elg�����(��2-j"�N	#S�*�U�9p�z�IQ���٥�?�]m��_�n����=p�D(T�R\�^]������!3w_r.�~FPO5���$�O< ��^��jb����&]vZvfh���[F�ķ$�&��-9�ل�Ê҇�n�������rʳ�fǯ�iט4����nB_k�e�[�Kd�I��xj���S���i@�?j�կ�j�GFV��=�g=�����<ҚI����]5�U9Ē�f���{��hxR� 6��UJ������Ӂ)^É�K�������:�W��J���[Z�����#O�+(�������5ѫ�jL���sV�x�a�JY!;����e�ɔ0��ʖ8�+ڹSW�ؿ����8%=��'\~d��e��bnU�^3;�LT�̐f��Ղ�8k��pأ�y�%�z{���-P� d(�!�
_�E��
���H���(z��HM%���;>+���8 ��ÃrDGV5��yB��� �r��G55�C		���a�pu�*]BkJ1�g���Jc���*�,jX�}:+�L��2�g����$N�j�'������V�RM���$&����V��'�w�Ξ���(��QFu��c �DAi�د�/��F�	g;�����3��_t��҆��yK����'�r*T����\4bx1������P��s�$ >�ʳ&��I�"��Q��F��&ؤ��r r{p��10w�K�"� �vD	�NM\F�l�},�r7�rr�-�̐W1��}W��Q���m�w���Țd�PH��tu��[��cUm[@x�1M8��4\m��U�ǅ�ª5Ie�,raiZ�x���Q���(�-C����W��	,�+�F��Vh0ZuN��~�5��mQ�G�Х����RR�-��T���e���(CZ'�܏��C�>��`�T00���H�,0qru���+���ȕsz�V�u�/��Ĉn��ۮ���0C�u'���J��� ^��q������Վ|հ,*l��w��[=*���9�P|9>t!2˷�`�|��f��D4��i�J퀨M8"Ƞ���8��.om��}l�o�0�Jq�����M!QB�A-:갨n,{��m�FG6C���ThZ�V�.̙-!UN��a�	���9��Et(LQ�\Os3�&�8��V�}Rw��IZ��yb�J����еWY"�-���~��c��F ��kI*�-�ȈY��}K�1�604+]9UL!��+3^6��((��	e�(T�'�RRv��#�7{����]hk�"O���'ˎ.�A����TY2�V�R/�p˧B��(��P(�3��:h&�
'>�U��Q��#B���sj�U�����q�4C��;e�d��y���$n�;�D?���<�����K��`�������y@�����Av�.�`𪱹y&b�)҂?T��U$��:�ݶr�4�]����ɪ�m�_P��;��@��ɾ^�;Ts͵I��6�\�2�G�:��^~'�����UM���v�q���f�0+Bd�ch����F�'�o^���6�Z�;>t���a��!Y�[2bp)����R��U�U�`��nC�;�k��4ԦX����)b@�"�>N�֋�K�hpj���ꀇ	J|�sS$ǟݯ_"���^���Z�ؑ)9���%�z���t�s�I�dWf�K��=������^]��1nwA�K{�k\^�ta}��8��Y���+R��On�>w6ꔴj��_�h!�����O�hV��T�Fh��+7"��Lb�JYHWя��|",��axa�������(ww;|���D�4�OKe�e��]}�ЈI��A���.�������R�;�9)�pӦ� ��X�@_�)�C�`�������v�QmK}y�2[b�p��������<oOBo|LniᕚC��ȏ��x�|��9F9��X������x��:�=w⬣հ�[/O4��E��e�p�&��#���G�..y?��j��;��ؐ��=8������(��:�C,��{������^�_&�ǈH�1p�ב�4�(q�Z�k�Cm�������7�D`b,��5�h�"�O�i�`��ec���]"m䛨=�k��9E�^a���l�F���":i	pqQC[W�T��Ҏp�� Sҡpo�t��r��5���D�Vt�/5�����#gm��b�=���{���*��l�C��!�R�����'�m*Z���j�2+�6�z9�S�J��*97�����q��So�P��UĖ��S᎓��G§��h�Zbe�7����.c�?ߴt�Tt��	s��Ai���N����S��������vK�Ly�y�L9\�
�ʥf�7��Բ����"�3;�p�z�g�>�R���֓������O��F@��3k�M��ūw�(o80�F�pυG�
���A��<<(}D/�}`j
c���4[�|{r�Q6'������z��ܞ2n� ��j��'�Q��RF�z���枷�u�'q)����A���8v%�g�B��/�C���JN�ut�W�`Ku��ub6�_Iv�H�O����"2����}y��az&�yقƤ]S6-g��˭[	�,�GW�w.W�L����N���,
0�q�=�N�dM�Xݤ˛%e%K��?{g@���ܝ�j�)��y���߫6l��ccQӜ�����edm���s�֤|��S��+�t��z���n��5q�Yx�IV�����[�+����XM�j�`,Iҹ������l��٥n_�!ޔ p�Y�O��R�+�W��7Ξ.{~�����)�������\�G�b��j0A ��Р���3��^�z�z����"8�卫[4�ٺ�
�X�T}���`{�pgM����%���y	�.�Ej�\Uòd��28�W�BFAA���
#��H���}��$*�0:p��'D#
�ۀ�n	M\�'z3��P�f��+�!��{AI���%"R*ދ4�E@��'&��ȚGn����J@��Uh\b��U��u20�]p,�m�(h[�	�7��m{��������|{���7l^�5��7�/��	�T��CQa��A����|�
�_w�FΊ��1��򭙿�[�3~NSu� [�����������43�0������:r ��jơ�T�Mڣ���x@�QF���ؕ��o[�T���UXW��ÔI��y�R��)��E�ƕ��Z�p%�)�ݰ����y���Ms�#=��E<m�Ђ��������{M#��;#)�U~[���h�d��������kWG̐���#WU��%*Z�f��[����X<4�#Xϳ�Kp��aB���p��?�ũy�������-�Q�7v���ܴ�]1�B$G�~}��z�=w�����S&V)ٵp��Љ"Fk8�\(���,P���@��d"#[��r$��}y=㼍o�ph9\�~_�<V�j��\��s�r�srH{+翾�į~lx��\�8��Z[ .��@��ס��N❆��d<5Q�'6S-�E�ӅF>D>��,�|c�L.���2��|����Uj��jT9s�]���18=37W�]�)�$����	>2Q�c�2�#S/O�!�x/-� /%����,��uc��T�P%So�8^��e��(P�S��Q�[chq���{�������U-C��O���1[4��?�Va,��0��z��h�1��������M#�����G�5-�x�J�f�\ �e����1/*])��T���U\"�L��{x��P��.�fyw������r_�BEK�^�G8ʡ`����\�JO��-�H4";# $�qG���)��A�XO�@c���b���f�3�VlS�&�NN�$y;2yϧ0n�
:��8j���j���FF��G+ @�� ��X�\�R��P�'�:���N�b��S��6�Q�R-<C�9Qmz<��9)����)�2������yˢx����i2��F�����`7J�:b"��<F�MӔ����G��-���j�o�5�R���4�rk$�����m�9���E�Ba�$b ��^�g�#`'2+|���#���
�o\3@o����f7E��N�="��
ZW���	VQH�]Vp��-�|K#T���xA
x��L:&bd�^K�Ρ�o |�)#j5���'�����gV���� �*��N����)�0G7cצR�1�bQ�`t(t��1�0��`I
�"GC'@()�3�͎�FfF��M��'�7:WW�Q�,��Co��lkBc���7�(v�Y{�mrzY���R�aND�d�Ə#_���I�;��}�}��NWC��318�u�?l�Y���k�啯[�����a^_O�}� �-�;�2L9�Z� �S�N\�*��r�j��qN'P��䙪����%tw����X��E;tg��
�Q>}];���1%mm$�=�,�M[MZ�����^�S��?��j�5� ͒�i���k�9?[��nFZp2�f�b�n����U/Cz5ǟ��K��_I"e,�4�i�ISeё�q���`�M*x���JQ��M=T�r!U�C�It⾨n� ���!a=�����I�xG��y�rV��Z���N	2)��y켿�t�%����3��{�DL�{�Aƭ�?����[,C%�ʼH4Y9���@!))i���4'og)=W�9Q?!6�B4y�ę2ߤ��e���N8�1�	�����Č��g���u����+��M���s�E�q0���;��R_,��d�D�_�DK���2�����)��]�~̨��z{�@�G�䡳~�:]������0�ô�E=ws�骸�i85:� ���EÄtK]��Xk"��?��JR��g -lQv�����<�j��<M�bc�5��[�[�d����%��n�������	��KTd������$�zZ�+.�j��;qؖ?�1=��Sd��9���	���e3��Vص q�o��^�Ax��?
{�ɾE��dX���sN�� S�#�	��|��o�������IC�������YL6��~�w$�߿��R�m�5��;J�͍�NkCx�����8�6��'(��~���ا5'-ȡKɐ��|��S)�'T@@<<����XT�z���6��4���+鉃U+��=�M�.�:�.%�m	zEit�0w��2�HD@'����Κ\�$}�������@��?(]4ثy?pUU�����8#v���%�[Y��u䎦�(Wj Q*��n̝J�v:xu�٫ C��< 
�F_���ί������u}�,�w���O7ԭJp@T���w���ِ��㟍O�]�5ܠ��6L�9�N�e����9�iWM] i�(YX0��a��d��ޟ��t���Ur(Ww$k����th��������$�F�����S�%Oa�!�S@��"�ǧ��q���"�� 0+�$��6����X3#$(;Qo��O�>��`�T�lSpk�|]�j.�_6�BL��O�,���h���������u��m�\��6��O��9���7���LL����6���� z��P6��4&]K�(,�.������W��6����#���8���s,Q�T�^S�W*ⴑ�j& �Z�Xq�
�/)]��/[*RP��4gc��\��<������/��a�aA��٫g��>%��K"׆ohS~y�٧>��YZާO�	�����Z*5�~������#�����mp@.��0UVؘ����/_#�������
�8+/Cl��8UK��	�WtJT9�m%zɨre���u��^һ��)vggK���%��{�73�k���s����5)�w�2b呍���$��X��6�v:�c����a��aՆ�e��TI�d@1�Pì����%X/r��^՘Zm�_)��{�zCW��G�^W�RC<��sL����Mϲ�.�н��i�UO#�R��q�a�7�f��ѯ�@�_i�� �����K����L4S죤�[�T,T�ZI�~� �Y�| .�O�+�e��q��7����/Ð��&�U�L	b��#��3�&��h�M �7|{ g,���rhƼl9�G�v��3�+�j�a?�*8�$�q�r>vA/���z#O�@Σ��. XGQv�-�y����1F�>��2��_ś(�UEqG�9�7w�_4aԯ�R����xWuO�Ե�a儤�KGӚ8�e��E��\H^BN��VD�J��oJz�on]���l�&l����P�o�-��>m��f�WZ������%G
/�ላ��mj��3.�k&}2��X�@ g)	���M#����K�����VZBp������?+'��U����T0ֻ�x�`C*�����ky5���q-jX�\�,�zl:eVy����̓6M"���u$�� �І¸(��Ǹ���	e���6N�gU�fkO�4�#\X�2'��齀|�jq��I�t�	ȯ�<C��*<Z8����5jhp���C�r*��kS�Ñ�81$��h���.`��ܽ������K�W�p����w^סa��$6��գ�Y��0������[�@~�"�[���B�'q돳�����.�Uz�zL��'�d(�,�c�,�U~x�2�EE(V�e�te\m�/~0^�&�?�Ũ��3s���a��]��c	CFYZOmG>v��>��
��?	j3˔J�}6�Xw��ٜLaZ�*�0�a�B/�iV�7�!� Ԇ�hS^� p뉲6&�ߺ_��`>ˉo����(w��	��`Ν/�욼=YD,{�/أӰ��5��Զ�⠔�>7c�)�lтm�B�J ,,[S���If����s��:���2nOT�\��#��Om��0��5-j�Z��d⣾f{Ո���N�pA�z����:_��v�W�Y�bq(n���@\���Q��'r�j}J�VXר$��>�ФZ���g�����-Cj�W�R�$m8��m�4y�r�7.j�^D>��4�h�^tng�s=�>�*-���BXz��dc������Wj6?.`>{��W�F9jL��s���pnuz��}�e����Z=���kE�w��y�0a$*Ċ:�Ug��XrU���.���U`�[B	�"�����v�wѧ Z�����g/R9��Y�~�]5Ac�jih��Sq��VTtq�_D0
��T����¾��Yq��瓝��~��m/I���Mp��$f������v�n�hD-���u���䵒�0]�H�#:ʥ�Bw=
�����5{^��� �#���m�G���4��0nq-�G�\e#'�u����Y��z���="�2|яW���-��k��$�T�,�ş�8̜�&��q�#2�b-<�<b`p�U到h�m�X�Ea�~@_��1������v;��NE�AUǠx�o�S�x�]�銇d�=;I�b�����?]���g7#֢[�2��9�d���!}��%�^�L���
��X<��=\�t�x�o����p8�en�%=+�6�����s����S��(��<Bnz�i��?�������t�ĵ�e4nVm�n�k���Y��*��N�%��d�Z'�VD�@TVtDJD!�=4����M�~/����O77�D��0����eT�W#�A�N��O��#�f0.�_i�h�,��CP�x�T���8�Faqvg(I��N�jbTH�by(~3�(h��?�xi�:�?�/��)����r�8��!9�����.�OiM�4��]!��l��1���~��U_ߩ�bR���
V�`N�
�v�W���i�H9|�qb�zAT�0ޏ�
�d`DD�o�j�\�)��Y��]�XA�pA-��t�ӓ���3��-�j�Iz�P�p�r�2�E�<������y�7 /`S��dj���� o�4�`�)��חF��v�,� �n�%��̼��V�S��^A�Y�a�E0+N�SЎ=�z�$Pu�T��4�� 4�RR����N|�9!�	�( q��8�Q^#:�yM
JG/R���������3��e�XS���lK��4������x罽��m�M�^\`R� \�i�r>�1��l3�t��_)�5�eK׺��|�Ot�?�E�IՀ�|�˓�����$��o�����r�iZu�(�JIޟ3��Oj!u�1�//اyD���G�G�^��D$��# ��}�p܀�}�re#��iV��o1�)����AXh#lH�؆��㲶�%Ә{�p�R�ǄG�#��K-��39<��̈Ǎ!d�����0��A�p�%)�	�Q����"�s��׹"	�K�q�`�"�g��Uw�\��al�G��+fZ��ތv��O
 ����o���Y��Qv��[�2ѣN�g�e:Q�6���\�T��F��J�a��Z� -՝��n	����F��a��4��P�ɕ#��B�֏)D+c^�U��v�a,���;�7@�}�>}��{5�oc�W2�1i*k��ӵ���h/�	����Aa_��]T
0"�ƍ�:���^O��C�q� Uz���W 5Д� �D"-)��k��q:��A��I��b;�5�������=C��6�'�X�����O���8D�����K�tix*>������?����NrD9HsŪ�z{�J/+�.��3ش����+��0X�Aq2e��R����
��]���Y#�	�����<�wCh�_�EE��t��L�$�W�޺���_��3i㚆[c��e���O�l����y�y>�W3tM:q6M�����_��1T�`I~���$��7
b�Ygt?9튳�����:T% ���@-�澥��ʭ��/_���:y���#^r�J?ۙ;�t��=z��C@��K�&]C�0a���d���D��)����~7; �����{a�ĳ{���+ϭ0!�@o���`xx�q�~/T�mM��W�z�F�h�f��H��TO�E�,t�bv���L�������U'����S!�o-������s#n�dI]�˶л�˄c �ZfH�g>׈F�۳�$3���n�5ތ�9��25���go��h&�������M`rm�+����қh�0*Z����d���;r��w�I�H A�����XTi�W���2�~�* 5Q ���Q<�v��蚐��{�����{(n7���"򺿝񽓾�����1]�a'��D�hi��Z�o���,���t��Ky�E�G^��ɥ�8�s��`J8`�;�3_*�/�Z�#����/��*��.u���Wb��Kj�ݨ��W���œ�~&O�Ș��e��$�%,�4|�'�Ua�W���V{9��l�o��߯��F�	us7CN!G,�ba��]T�-eI�w��>�z��c^�5���N��[��qh�Ұ��Az	o�$���������u����BlщX�M*���NB��:�������ӝ������s L(�ɥD� Q��^ۡ�դ�ӳW(�F��|��<��3�YAKJE.����8�2��tB��+?���g�,� X� L�%�;�f R��^d�\ ��5�2��L��ْP.x��nI�O<1S���v� ����t����.��<\�F�{��D$�ئ�[�k8���� '�S����By�Z�3��C)o3+~^#�,���>���\��<�w0�#Y�{�ß��YU�UjU�c�4�Ba���i+eGΟ�~�EWl7|����F#�z �A�[ �v&�2;=�Iiņ��eXG�89UAw5.�$ݦ,y1��'�	hDg7���c�#_t�a�F��I`��KBD�e���~�z�u��1;-���x�T�'����N�|��]��f\\l��m:pQ�Q`2�0�p��c��K)�4��)%�� _Lg�� �{]0�y���eJR:�ߴ���55�iSY�?��hy��h��ĕX[�0Ѣ����/A?���l3��~$<�}Ƀ�N7[L�e��Ȋ�^٤�[�<�;c�/��
��I��>�y�I'>l)3|�j���E;v#�ᢌ����r_ewp�09���o�#Ŵ�8t� ��2�v��A��N��{߳m��c� ?��1���9p�!ܦ>Ш���|qtI��������V������ᓭ���Z���)r�W�	C��[�beMH��J�]�����g�,��	 ��bFt�O'S^�&�Z����-��m�i���H<��\&��d�ߵ��2Y�R�DR���e���7�{jW0t��d�yY��q�ZO=�^�K�.��u�U��{�}����b���Fv�c`ӹ���:fXk�����4ݫ�v�;iVL�������aD�����Q�gI�}���6�X�K�U)h�>!A��Uq��ϯ.�ux
v�j�&��P��ow�gr]o�w�N �ZQ��Rq�
�v��'0���yxL�.�p �4*����?J;:!��H�X���5�K2���]X�N�Î�ȍ�{rvni��Lf��%_�-�Rg'�.��������s܆�o�`X+ŏst��D����W���"��E��c���H�חmq[&h��X�	����ޗ�� ��O;�Կ��\��#�F$6�C⒉�!�A`�_�Bw�� �_��f�8��u�v1jU_�-�LS�
?)K�N/�Q��%a�a>Z2�q�r����i�ӗ�)K�M�$��茒����$1�c*	#p�`�K|�z�>'�	K=*�\x�`�Z5l&�Sh�Z�ҕ�G?���9Q"0�L�2Ƒ�VG�f�N���
�����9��%�����'��[)��:�C�!�*��=g~���Iy������`��8Ҟ+j�,Br����%]M�A'۩naa�&�F�b�Fd�dH�#"*m)Ͽ�g:k� V<BB��Q�S�	@�V��C�_�e��d01�5��?�t�U��s��ԃ<�7 ��F�~�I��W>[���i�G�,߀���/���w?r'�6[B�ۛ��,d����$J�N@j���9�f8rښaY�T�:���F���;;�z�e���0� ��;(p��׼��E�_�	J �UQ�!�������,-I~sp�����1�>O�[��gw�YW"ހJ�A��]+�`'
*��L���"� u��p�RX��D���u���)f�Y+��6i�b=Լ�9A��>���WPo�_��SLf�$�z�J�Ә�>�N���C+� ��糣��tCoj�d��F
B��3��	�.vvYt�W��$�P�(Wh�cjT�ć����zL��,4`�5��V�}�[}�4�K�V���VP�$�tgt�G�=�J`�*�};G5b��#�GW���ĭj�]`�ޮH ��-����-[Z����k*������q�$ahH�$k�jL�jacc*�J�#B�k�.�<I� �O����$kP�E�̱ȳ�15�����i��B������G���
���*�Z'�wZ9@1�����#���͗�<(���~7����s&��~�uL-z�Ѩ���n"�W�\��=�}����[�{A�Ւ���fm.��/v�̹T\�i*��/W�� [E���T^�����\*��mJM��JA#��"9���CNS����Z_��3�U�o2D�G�;@TdR�@O��mA����j���ʜh)�	��&��x�ƶ��v�	k3I�Rín��g��X���2���w'�o1����b�Lxs�`lg��6vq�n���Q�UG2��\gB�Yu��h���Z���l1TL��"�^�m�zT
��J�LE���57�Z����L��}�0���AS|�VG���0������a��=�ul�c
!-/oH�\�n�������k����Kh���2>^z������`�^&����J�	�	X���q� 2(�����Ʌ'_�*����[o�cx�K��'W�B�M���4SI��Z��f��=�>�^���S���z��ea�
�5�ߗ��-=���^\�/D~��ĸ�x���K�9��~K#k��N�Q+�MJ��$7*�b����l�G����#�D��t���żP_�<Z1�S�8R���{>8X�M�Ǽ��<���Lz=,�{�5W\�F:�n�4�al�,#o|���2aY>�g��val����l�ѳ�&+���`�w��� �f���B�Em�mX�4_�!=?�`��-�����6?U�+����ϟZ�	�_�;��K<�A��5/R��|��qs �ص�
`�������I��{`�Ȉ���kQ�����ߤ�6tx��#�+x�SaE�h��{x�0
��6XR���,���_�n�"Є�]^C��o�X�;Ҹ���Q2�7��\P��NJ���5w]�2�>ů���ƭ����Ӓ�vl[;���$)c��Q�������!I���~5䷵����E�nt$e�[`<=���5	���+:VY�@����Ţ�,>�`�t�`��eH+[-���G{��ko�i��s�C\����w�,�U�8<٬���zeo�+�ҵP�.���_í�Vw��)I�̜cGkd"��ަ�"����.>��6�; �C]s}K��xT����>��V1��B�5�J���%M���4�����@��ՙ\~6�n�Vx�c���☿�%S�;v�;L�<����Es1��\���6G'��)#�P��fk�t�>���;,jjvEVK&�y���(r��b�^kzup}���W �19�ˑ��mV��s�j�lu�s���-\B.��#�^/"�SǴN��5�����7gVn$#OF����}܎KĎ��b:4x��X���?���YN f-� ��xy���Q�!;.����^����]������e�狽�P���q����M�9�T��#�آK��g��Ց%V�t����������Z�?��d�S��p&�"L
�>߻�� ~��ܜhI�b����/:y}���p��<g罈��
T�0en�i�a!e���J�Ra�q�J ���P���r�&�l��-��/��\����o�wn���lk�N�d얄�пn��v��I+��Lg��ZL��n�Pe Z`�h]�Ғ���Y�zo��ndF��-!9@��X^�śY��w�H|�Cu�S��
I	�\�:��B1ĵ6mλ���P��Ϊ��_�3�k@tb�XR�g@�k2w���.�.���t$����㏬lӣ9����3hZ'�
=Q۸�X��� ^�?�h%8 �D@.p2�(�PЊ����.��qT�ek�)Ɠ��O��dj�b������*��z���#��-ͅ��e�4�����N0U���k������[6�>���]bR<ٲ�Y#F��U�?G@_1�l���U���N�Q)⨸�R���a{���,$@���c���rk%�FV.���Ǜb��7
>�^��|�o;��D H�SL�`�����X;���E$[��5�'�Q��O$2}������q���I_K>;��*��5�t�ؠ"'�d!�e�hu ^�:4��нZ����X���B���R��>����q�bq�Pώ���L�ᡈ�RL����=�n;edfj�Y�*9�'&��{�%2&�33X�3�;d �a�*"zcR�	�X�Sf*|���\�t�C���袧��uGt��J�8��Z*l�V���[��0��y�/{���]OM��$�9]�]�<N{���g��\�l�e=�S1�����!k2�~�.���(,��FA���d�Ĳ����Q[�,��#�j�Ln^�FwM��*�)������Ǟ �	��1���l?E�[���z��z����[��"���e&��>Ŋ|&�a��;��Y�D�1p��Q��"��PG�m�ɦ�߯�1�������FfqX���Kr���yMHDf���|�|&�0
�My��Q5�e)3H&��[�~9��	���ҿBd4���/*k�-TE��TM�AQ��"��GMʬ@**]��,g�ŋ1����E���o�X��x=�z��3��#��Q�^�F�m��V6�U��s��'L�ι�]���m����d=y�7hZ�0�����}5F�%-�����iٟ��]����Q!�9�m��'�6��?��)n���`��S�xŔ�h�zq� �殞����DE�%�s��7�rƪܛۯ�5>N77 ��7j!o�����lޣ]����1!:"�jl8�H��ƿ��nzS�5�w��Q��b%�BM��d��d��&�<O�6�00Pt����S*���U�w��5����Ǣ\ ��:~Bru9���̺cUD�>�!�d��v+�^�s��0y��y�J��!���
k�Gbn��?��2��&Z�-����wwww)w�ॸwwJq����^�%-��~���W�k'�f=�g�d�+Zx�����<�F4K�{�F�P<b�	�TJ���4�T�`0]I�u�I�DL��.���5�\��5��A<!�<F>	���I�_�5�������h,hhH2dɰ����MU+.��'1��J�'&'ٲ2��6 ���bT!J�l��0�x?L?E���$�2t�Q=���v�@=#�Y��h#1�տ�[{��oHBC�ߕ����(�G������f�]���}�ŭ�(]� �c� �������NJ��w�>��n�3ty@ ��b�]�����(b '�^"&��Jb�X��;P�"7��MԠE��V�5~z){��{��sr3��5�g�s���H{��ËH��d�&D���B�34m>C^���]7�])�O�?B�[��ZR�����6��/T����a��Α3�{�4�|)�*�Y�j�"S"A�O
_���5`_�7�K�|�����b���<5��?�#4Z1-Կ�86p��8�emgc��;r����e��ᢎ��H%����_�g���eyې��� �6"u.[vn$6�6�h�?Q}D���+�1��nRT�9�����ЧAD��*��OXN� #�<M���j�9>��C��+����2�S�M_��</[��I�<ѣh#Zh��́� �G@�
�+�����)7�ƾsг���n0:����hD��T�1��d�0��!����p���1}�W@X���Vk��S
K�Y~.����^����l��[Dߑ���~�J�%q$YZ��w¢b8���&��I�� ��fe���0e��K�8��4a2C��Y@^I*���"P;�����u ���Q�
��]燌����Z�|WU��M@B5"��i�7ά�Ʋ{�$�t�V�B��juZ��C�r�'��<~S&ZS�Q��Q�\d��܅'�u9<<\i�b�7���)� ���{��I2��4(��a��s!]��w��@�Be�YU�}B�W�e㟔��q�y�R۔���"4e� N}y{̨�H�B��2]z6.!��O�
�G4r��ysu���.��!!��A]Y�_�<`v�%N�0�l�x��1t��������뉠{wO{@{%9#�woq��죶$���!�L�|���.�X�a�DU�A�,ٮ�l������]��}(b���G��7k��C;�W��"(Y$,��A� G���I����=�������7��\f~Xm�<�'������d�j����P�b���\�n~QgJ���R������[H>��9Vͥw҉{�;
�-����	Gk��m7T�E���I�s�~�������U
�vW��/P%��TK���Q?:L�搣����?c5:l֮C���/c%��NV���B)��A��$
z��|������=^�*��~<��9
��kAT�,���(��im�n������g �4U���t�$UWf��������+H��	UG�ƃ�X�;�J�{�����/����P�2�P�C-U��@
.�N0,\F���K�^�V����S)���>o�O���X'ꆊJC?f^kVP
�����;6������������e���Y�5���Ig�g���0PLU %]���8�,9z,�������
�>���~%F�!���0~;�� ����F�L�p�ͺMrܼ�I;��7D��~]|k��A�Ʋ>�(�\��г���+[�k�!�/s���`pI�P���x0R��H�;��հ
�UN�s1D�+m��`̏ ��;�u���.��#CZ��зԔ/"]�v��)�A�$�q����&�e"nG����{���!i;��Hڼ���W"A`�3o��5��߿R�!���+K�Jr��ΈS�@Hǒ��yo<f��b��a|;
����L�Sߺөvh�aM�q��*Zf�z�A2��*�B���$͛��8�	gfI� ��$��;5
l��=>Qu)�$0!8��Mʚ�w=���a�x�N���r*�K�N�/Ɖ��L�e�֛��D�/����صV$��mP�0���G2<��d_�4N(OF$�i�Ȅ;fŹ�T2����.��H>���Ҽ�,d���e0��aS������Dh���5�B�rrn��W"���cJ~���������Z��d����a�Q蝱�J���*��M������� �{��)����������-c`�C�3~�6#"%)�����t1/�7�[`�Y����e�HX�~=���V�bh�)��:��z;y����e+��t�(B��������1��y�y~e6��_Y���NV��.H.Ԯ�]Z���q�Gd��;��?11����t�Ka)hP�� �6]6������Ur����ޑH*(i�ݭ��z�"���i�k�Q}�g��})�����x�\�ݠ�??"��Ս��&�inٹ���+ͺ���V' r|�ר�(M���_�.$*�g��_ې��2;���\��fCxF�~VCx:���J�d7k��m,	y^FY[U�����>�<��x6�t)��h!:�'}�J�ٸ�+S�Q��NN��T��
��ZK�h�jMU������U������>��
&�Ֆ�%U��!�(��uDY��r��[�[Bg��e*�ݞC[k�+d�V��R���͍ۓ%6�<�F����-�������-�8�����U�q�@�n�[w��Yc���%��
]�L��q=!ם��v�l�[F[�V/"�愶n��]v���q�S��O��9�P��w2_V�ͰpƜ��BQI���j�Ÿv�$%���T3�A;�w��X���ٹ���9#�-r�7��8F�XLO	<�B��q�����<[֊Z�����
~-O=�Թ�n��H��H��<��P7�iF-#���X����%�Ӈ{����ى�U�T�`�X��@�Ce�p��\o5�]סƦ�CJ��y&���J�ކE�����)6����h�p<-��,��ա�G5�hP�F���#�*���w�	
���bp�c/R�=(�L�T��d�R�P�j��0���iI���WQ�Ur�X�ϱ���O��z�	ӕ- X��7�R�5��Jv�<nn6c�����V�ՠ�5�ۄq^�[@ў�h�k��������lA����bz�f���/��]���2auBi�
mȣ�C���H�ڨ���Y�Mp���Nˉ-<:�Iǻ���������� f�qwxT.,,x��h�#���b��U[Z�ݲ������{lfPb
.�z8���6Ҭ]�{/�9GP0F�[��UHm5�ަ�ڮ'z'�=m��瞫Q?��a��Q<Ĝ"�LPy%��ME;����m�ۇT��u7Xo/���\�;�~4��u����Ju[����{�b3��呃z����u�˿��/*�Ot�|�B���L)��Ϝ�!^�f�>$���ZjsR�	�C���R��_����cnp�͍	��%�<N$}e/̞��М�e���� HV�>�[���hS�"p9�N3SU�p=5S���H����S�S�o�&�ߊ��c�8�0�����H	��5�
ϒ�3�\΄�|�w���'�ڹ�i�e�m'-�S,l��O8�K-R��
�ԭ?��͂	f4�lll�۰o��"䃚k'���7Z,�aay��Q��Aˁ��t��o]8W��V��U/{"�����׶$�-��l��3��D�1�m�nn����_�|rT� ��?���{��z�!��c=��*$Q����������EN�>����yӏ��
Uy��������RM:�Ȱ�:;Z㧱�z�ef�;�d�6��������x���1�w��r�\�"

 �5�(Aす9%#6�^>H�]0A��X��q��{��\���#F���"*�ٴ��Y5o�tt�	��m�H�j]|RY�/ ���D��� n�&�f�F�����s��q��@��'?x����r ��WUΡ������~°�,jٔ�Ў�L�fǮ�]O92��ʴX���� U���Y�����\����E��RZ|�Z����919�S�/��枮!������/�]�7�з��ֻ�QJԱ��Oڰ^__�{�P%��j�_�[[�m?����J}M�EB3����V5���s���5���q��oO�ܽ������v�l�)�YՐ��V_���,��ɦ�b�`wS0^�H�t�GBBBQ1N�b�����{7I�ze/���l��-QP��y~��~�lV.�Y�͚K�7��D�;��(�Wʬ\a�ڭ")� ��ܔ�y�K�z�w��,�f�z�$F�������N�`Y���9TTS%PK���hP�~�y�,oe����:gj��?�.w4�Z�t#l��<S�i_8����?>���%�;�?X�hsx��@\��	�!�l����n�L�#�c�CU&�1k�Č�|:�ԫ�Ȭ����BV�I��WL#:/+�;� ث���*B��i����i�R}���`�0��g>�/��F.3� l�G�@|S��a3�1~�.u}ْ����V�o3�bjn[E��F(??�a>ޏ��/XN^�/�?M��	���똲���Ĭ�b�T+���I���=��~{����znJ�&�����eg�p�v�ݵ��-Z���B+CO7_���� 0��}gV6��Dr���s��*��A�M
��# ��X���OPݷ'2�pb��e�X+I��\����q��D��4�r����0p��pL랄�w�,C�H.e�Z *΃N�b� U����r{_S\�[���p�_&���W�kS8J��	�,1
�7Y��!���C]�0�@;��c���[%���i�廇�p@����G���y�]]T�?��־��GrT�|fccC�#�߮����&��Q���f����MM��TI��xf�M�v ,�m�"�Bn�5��7���4>�8s� �P�(3{n5�- ���
=3;���Xs�'�4{����Q�?��OTq˭��'$��WG8�7�+��y\w4W5g��z��6y�񇆅��<g �k�.o�"5�f�u&�f�rw�#���%Om����=�`6/�$"W��\��6~֤�f4�ݘSlҧΚd��Mx�e�r�b���*�tx|IZ��v�B�9�8`�{�qnN������e��Q�,�	������܉U���+@ԇ���4�`z@���;[�6w��F���]������X��a��]K�,�vUiQKx�*ߖ �؊a�f�4��W�mWVO8c��q�D�J��0����BU:7�c$X���4�������@W2P� 4��M�Ϛ~�H3
@�VHN�e�@��~^^\
<+1y<p��l$�YK��V>��5�'	�(���[T$ѳkk��Ⲍ�#��G�Q�MS����������kt8Q�Z����4�l:��e�i/������[y�^ˏq�W�����ι.���#ۉ>����vl��
�C�'�~�~��"GE�L�a�n��7]�K�^�x-�k���Ҳ�K���-K�?1K9/��M����J�DR�v]�W��+Q�YJ��b"�`g��|3���P���R��	�|=�,jo
�,���4s	�O�.-+������T���~��v�"�/������5��!ۇM��'F��k���އ�|��\�$��ME��;��Q����xd�vKH��&BH����cX[܈>'�o"hRP���e���v,5d�|2����,�-|�������r�x���>�ļ��@���H����K��~i�6�c�X�?�F��0)���~����g��r�3��.�kq$�rؐ���3�ŪUk���2
��"�/	� Ap�3���~�v�G�Cg��n�]���]*�n�<.6~�]3"�}�g���k+��H��wf���Z����ͥZǐ9������:��E���(R939r�Sm�~�b�f��V��b�eM%����㌧BȞ���� )�f�|���H����B�]u��0E�w0ȳ�ۖw�Sⅺ��a�)��:'�xVh�����k".���RDM=���׌͍R���6Y�lɷ�cǴ����&0~��t��U��ѱ�~�p;���)��*xsh�B$ ���r�5����؋�?�����S�sn�%�vHN\���@�� ��dI�M�s%ur�6=7s©��hϊC��8`�3E�E"����g��o^���0�윗�MĀ�k�'�	�Q�����f�������%G5�=��Psv�&M��� �@����!ԯ]�7WUU�y=����C�(UQH?�������`X�+�ױ�~�o��1w'S��@�����>�C�ނ2��Ը��;���w0�r��u:�������~�%-i	�񇻣�,RN��R���*�Sn����C"0&h����=$僡"�G��*�if^��^c��ũR�I>77��P�ԛ��|?�����áɻ9�Ѓ����A����hj��;S|X&�b?i��ߒB)��8g U�A4�J���jC��� e��h݈��������$˜f <x{�4\1�җeőEGX�uoBI L*M�Ұ�`�ޞ(��	4�C�W���Kß�8Z~Ϗ+Р�Ca��t��LP�mB�4ըy���t��Cl|t����ot/b�����������Q5F�p��D��Vq�s0i�v�Zѩ슻fIiܽ�on:-Qz#��Y�<D��H��,rR;�������+��)�p`G�F�F����]����x%�B6���{��~�y:����o��K�+qA
�#�6ׂ�U\�{��}��fj�uTCxQ����OO�����v1Q���Ohw!� �k��y;�^*�L����T��m/c 7�+�E:��@��8#�}iP.�r��,Md�@��+
C�<��� �N^׆�ob�wu�þ�9��?Xv����2�����?�v�oѫOOfñM�����E^��=���A�I"�,kn�8�D�:Qy]��1�/�k)�n��Z��:#�<<2�i �ϲ� �b]2vt�_���t�x���������C��I�28�1D�vss�[���u��;��/�)�Dg��(�{~b�K�mpDp����>��\o����?�7���������7|���� ��(\_�A�S"#��7�!��:�����" �"{�[��{=x�ל��|��¦�.clo�&#;7�<#NQ[U�V���C	K��.G+i����!lс��XFE���r�.?9}3�N 8&�@XE�<���ŗ�'F�ԉK^������3�<	����Y�a�a����a��ȑ�;��0��(|�����=�����nE'k�y�?��f�'��m�0���ɰ�K���5��g�8��]�!�[X�Vr�k��=�yɓ_�����Q��H�
�2'�����M1̞Y�I����
Q���V\�G3�`�Y�/��W��a=���	�luBub#��'|�`v�֖�[�����9��<�0}� �������5 ��t��H�&�>�M�NW�Y�u�Uڴi�.ӗ���>>>�%����t�]�,��������	O�b`��������Q���i���<ƨ�cJA`���!'O��U�ocːc����7G\�瞇��A[Uo/O��F!�^������x_��u�k�Q�=����8	��--�\n����o��1KK�2�B0��V[]����9lb������2B ����E[/.��_�v��fff��8����Ld���*H��$Ge ����/a��4�VHH��u���W�}ܝy��w<�H����0�v���� ��J�$;'�6�fgݏA�\�V�r�7;��=��.��KY%���0o�[�A��^�0�k��?G���]�U�4q�9�`V�>��iyIb9+�D.w�=E�<��i#�'��$L��V�e�܀�r,+���\�i�zƏj��\"J�A�8c����=�����f���T�'��Z¯�*l\\R**�,�ԿK0ƽ�XMQGv�3'����u�C[7H}�q����/hz�"#��Gs�
C2��F~�ʼ��o����Z���6^�=���j �Ӻ���~��Q�Z���W�#i����L����Dq���,����p�o�]�[�2 ���J�����!����i��ƩPʴ>q� q���̸�y�S�QE6M����y��YyG�*BSN�C:�W��
�3�Z�}�g�%�hjJ)syk��X����JGy�羆��&�,�i������������Gr>_��yƫ�~p�r�	Wx"�2b����a0z~��\_*N��"{_E���Z��A�����	+^�G�E��>?�v�I��*��#�;�~	��I��bSقRnn>D��'�uO"�[�f�վ������>��=�q@�2��)gwz�&��H���?rX��Z���J���K��g�i?�#.�C����_���;�r[w���!V�8�_�^(n�v��FF~��˳���݉z�P�����I���b$ʀnC?ǵM�\�Ƙqo�B�.c|`�����a�zX����F����.)�PY�#ّ��31�U�b��?��F��p�S�~��$=R�.�!!/�$Y�d���/����*�	�<�m�w~-�5V�������sf^�E�w�{��Ӊ��0��m����%o��πb/�1W�!�2fH��i�����i����o����������e\	�l��X0_ec@y��1=sP����/k���JV���Ay�}�	E�!�k{j�N����½aכ�C�9����p�	μ!'ˇ�n��S^NNO���h�
ښB۹��= �!?�hc5��\��!5n��I��@F�Y��[�,[����N����@	�Iv��Ƿ��*��D�A����FAA�2RT�� 4c�P��#&��)��p�9A�/ ښ*���(���V�W[M(���)��8awvnb!��5�q����p�R���R��A��.��cm��7u�əB/x���%F�W��E��=u�����{z�1=��C��_�/�UD�ݾ�Amb�@����^��ְ������2G��������Iu���4D 3�̬㋋���,����Q�X���L`a�.cT	+	�ȷۿ�{���2J�t�h�	���B�ǳ��������3T��p@���\9�|r{m!*�D�a׀(��Q��u�Fcg���7�=� ���Y��U�.��� q��7dO�����sѴ^M�@3xn�8�>�d��\�!3��e2%5�V�m��i����O)Ӽ5qA�]˲���T�!�+� ��Ư��1^��%�aey�͗�K����T��ӯ!^q$V4�Q�$k�G�G4^�����zph�+H~RJc0�܀gD���ux�$�F'8_�Q�υ}����v��£VyoR��a'�����9h��ʞ"��T��ٽa^��/gWKK�	;��9DG���u0�Hs��C:Q��F|��������/{x_͠��˷�cE'��I�qC)�u�ɧ|�z�t��6�Sh*+���B�=J�c�nz�h��C�3|�w y�?���Rlsgw8:nw!.1�9�r�R_��
6�����r�Ļ7zD�Dz��C@ X=�����O�d�c�0�S��j�^��p�Q��1[bǷQ����xIi�L{&I{���Q�iT���tjF����2��诽�\=�@���ޙ��\' ���I��յ)5�fWWG�'�`�����2�-M��1j���C ,� ��6�z"��B�g|���jd��p�?���z�ڐ�����R�Q���l�Yh t�,=�)S�8��<c�����ߎ�o'ߝ޿��C���X��c����/,�4�� T�I�*��r��-W��2��:�H�s6���K��©�#RP�Yedf�WP:赪�FK���6�Uq��g+��)Y�+�$I�-�� LLǨ)��`�YZ�D�-=��:�����FRt<�ux���Jr�m"�<��{�;�[&�JWdVdm�	�g��}���$�Y��f66~6b��	��$^0RQ���A:�P���p4UI�w�������vS�1l�]�'�_r�A��$���vw@&e���ջA�4x�c��#��x���m�k�E`�!�F���=�ඬ�W[<�,��ڤ��h�P`��cJ���䍨�OC�eTe�% [�LÍ�M�7�e�e%p�sLnnMXT㙾1%��8Z�\�ض��\�1CC�n�W ۅV�=���?��P���"E�8�e$b0�OvIn���C�K��1a$@bC[�qh :H0sQ�_��5�8	�ʖp 9����flPrHL��%&4tt���R�D�m����F.��%1���wz'�/;zj{��;��SXJ�*��Ӣ��g�mvY���T
�Db��lv�㐈3?��9.���pK��" E��a]�NiМ�H��du����Qw����Qɤ�^��(_�'XCOIi4`����ܵ�d�� �)�t�����J�ㅈ�)��f1�IF�i#,:Ƴ}�!����y^�fa{������ى�`����)�h���(���?ٷ�x0�d����3:�;�&)I��&>s�q�KbZ��KPL�&O�I�@�<BMRMe,ܘzA;p`��h`RO1�2����5n��0�x��.��6k�7l��J�w
���ո�t����NO6,�!2�#��%�!mw�-��us�\�bDt�6�_T�a�9O|��'i�#m��J���5�O�/E�мi�W���qx��l���T���~������s5���cӷ)�-���H�Ι�zϭBUY�γ����wM%m����
`c�S�E���u߷?+R�abl�P�E��(�k-3�Ud��p��F����헬~=��:�U��a��l�,��NR$�?>��� D���5�J��m�A�q�Z�4<�AR���w�Z�PB��TK�43�,J?�����r�j�Gw"�U��F�ޭ������0�a^{%�B/�$�f��С��v��R&����%�����<�հ�K�������o89Lu���8A�C�>7�V7�9���(\R"m=z�=���":���5����nj�"��t�m�>��p�u�m7�s�����U�9�0�Ԁ#���V���\V�d7�;Z�
H���M1M�U.E��?��E|In���Do���l�m��������vF������9��`7 U>�+7%vЏ���<bL|����=����$��yƥ����y[�1ꑡ��#i"GV��=@����X@
<o;2��I<�"��X��N�p�2IF��]��!��T)6H���g��0�p/m�2wqm�z�DdH�+�G�f�W(Nފ��&Ga��q1����b52���V�����Mqů��4]*׆�lQ��|�:y,%e�J�}��������4�*ea�����~]?��rf1�Hi�K��&�m��A�#�^����r|;>K/��d�(�2Ts?���Sڽt�}�4igp��y����ѹ<��qj�;F46> )PѐH�L�znږ��D��r�G����Ǐ���{�`�XK�wՉ��j��ߟo�/�%��g��j�Y8��M�S��>��1�e�i��bn�]��F�$�?��s��>���A��4V[��=x��tH�f� ��#�i�?ekp�w�d����ץ`q,j,���t�L!���mVB�F!���������xņ�J�cT���11����¤���2�i#ߕ�	����Zʙ0���_|/�U�^�s�*�2���������y��2'G8�n���?nZz�3ʲg��7[{�tgju�BV��7���N�8��rM�3>�Qv�����5s�&���j���"x ����|s�4��U�_	��m4���ȿn[,(k�ݭ�z˚T똽s�rʒ�� ��bO�p�n`�ܾ=�9�Io�.��w_���R��FU�j�穐�s����[X��79F}!{ �&����F���H뾇F\��AJ"΢�+=�h�!��ٗ�R,�)�J��5����_veKxTHu=��G�;��lC���c6�Θ����w�,\+R����Q��,�F_uJ���K�"�����<��P�]�~k���Xt0��4i4���&LZ�T"�浧l�a��]��
��d���æP�@<4�k)�J_��(�Ă�p��҈_�q����� ׿,�[�C^���+!eO`�j�E�N�LV����qT�31̬������5�:-�Pk5M�}4����²�,����#�Y�!nP@#Ά���˄�V�[,���p�8e)W��[�5}���zB4�}�IҐw�y��ANX_>��-?戼P.����~/��=���C����L�G�ڰg*��N򠆽���Ȓ��wo>	u#��ŕ#�+��,��!2�����љ�mZFCE%ζs1��Rid�x��T\/���Ɯ|*�];�Z��u["�uJa�f��G��異���8���Q��w�m�
�&Rlh�h>�����"���b��&��v~���b���QzYK�܂cҜp��D׉����ײ�I5G��gr�e)��%�!�����B=��׉�	��I���d>�ϟ�/}Pk'Ȏ@�;fJЕ"��;�8����7pz�r�$����=��Z����V2���I�\�z�&��/2������y���ۧ$}正vA�#�dV���z}2v�ݠ��^F?�/�MU�!K��rr8�2����b�������aދ{C�R��81]���Q^I��`lZ�H�o1_�E��:�#rV*��[~Pɰ�hѥh�m�z[Z�oyE��ں���f|�..�.8!3�U�R����s8n{zeJ�d�x˶�٨p�	}�[[�K5(�2��*R�; }x�l`�_C�U<�|� ���8�ҘWa��9�0���{��֚�.;'�,�"ҶSY8�6o=�}mɕ>�K`dB�!�o�,i\����<z QTR��E)Q�d�c���k�
U�s����>��u��k��$���喽�!#'s^�:���;�ʽ ��
��D�ګ�*�*_P��-����aA��ȨF��-I�A��!��H��!5i�,��8,B���=o��$��❳.�+���ْ����n�m�����g@,b	A��rur��D�!��n���n���	�¸���B�G�ءa������N��Q�����J9r�<�+�̲�ۤiڶ�7�,�/5���*,��������/����w�e��?�A�1�Z�Hrp=U�匣�#u��FP	V5B]I]����jF�ߩA�)A	�hD��=DJq���KZ:����e;~Vf����3�	濝���*l�nBYh�������!Dɴq�JZ�tN�z�������G�?$��4��F�-�TD&����n`�m�'�§ͰL����;��	+ �y�����tzۖ�����V�*�b\�-xf�)��^(�Dj�뼸����-�i�aP�k5k퍧G�{u�;a����8�[Ƿ���n=o��Ah�����%���#�{>m��lk��/i����"=�2>��U��N��f@"\��_�����U?�����h�������y��R&��h�V;�x$��sgMP.�h�
����䋠H�m��đm?��fue�`�c�	�O�>_�$�t*����Ũ�$���:4�̰�,������'�^�_���u0��e�̨�l&�� �O,9B�G�G.n�7EE��~�}0���$�=�l��i��E����7b�[��K�ǡ�iu��dBd�*�>��P*��f��z�_���d��$��)�"�+sd��k��w�ˑ�z��%ih��))�	I4�Y��o�9�Y��!�.&	�1��d�P��\�����l�	�����yԐ=���j!�gp��O@��a	����FR�٦Pz��2�x��^����Y~��w��^Q&yx_M|�	 �Wf숼�nI��z�R7�+�/�H'D�����i��+\�1=�H��U�]u{�+
G����x�:�Cl��z���6)�f�2Q.�Z��87�Ѧ�%����u��"�KVcY��B�o�)��	j�9�*9��T�>-{�̹�z�O[x����n��m��܆���6�֠O������Cv����g��j>UpO��k0��/}�,L��6`:�W|����u;�
-��eζ��I  �	��p�,^M��e��Ե�>�hU��m��#X�XR`P�H����`� 7'g�?t0
�������Y��K���E^e�eWYB��H�j�fdd]ٮ�-�H���ʗ�x�҈۽fm�~�
�kf�N<oF(���!��w���Ȑ'�w;m���hZ�0Yx�ϳ��1sd��ä����"#&}r�+���\�O��<����?��`��������n,s�/��p���J��O��d��00��d]�0�o�_Wk���I^�X���h#"�ԋ�#����)Qwa�����&�m� =^.և��d\��q~5�K���YF0����j�p�hW�U���8�'��w2U):8|�֓zȄ�v=_a��\?����o�Aŕ��"��.�2��hp+���	O'�|�Q[i�+���P+E���K?���L�:#��Ųa�����7����'��A���cs���'��%��mG-'s!�G��cL�����������w<Kww,:�.������5}�jVIk��f^O��Ѻ�v�%�4"D����b��5�8M�0��ԙS-f�N5�0�IL�>��rE&�U,������Ꞟ���R5q2T;��'�c�;��<�7M��M����BE�G��xz����Yp3�,<'�1�"�h��K..�ΰ�l���;���ޛo�͌�G�������2kڹY�b��	s�5�^v��l?�QܦFAJ��k�vX n�YO4�}��eE�B������4��3�&׽>Ȫ�8w���~�&m�!���SQiֱ������H.W6/KǢ��_�b���%_i�8�cy���q��qiq'q��j���	��n$����\��ܡ���������a�j~���7^�����&m�����
\O�|���X�NZZ���2��q�^s���+LF���J�e>��c�m]��E:�B������^���M����
AX��aщ(�&��L�v&�� �$4<�1v��A�s�p+��@{{�j�^g�D���D�xB�'������2|��Kc�#��`�01"�b��NL1o��ڛQ��x�`^�5P��P�E�e�hs}<,�;,���������7��!x�Έͣ�*e��XJ�J���+�U�4�k&M����0���ogt8�D�$+���/�r�C�����5XM�W,��Q���Ǝ�s���u/�62��\���6��hV$5��Y��p��#̏��fv�����V�غ�Sl���+��~ t90U���gX}[��.�1�%�`F�Q�k"�Cw�)���1o����m�6���Yᓐ�HH~�9d'�<b-¤��wT]])^�51�i6�nJL�:����s8��fB�25g�T�y�6YW��&,��z�!N�E�B�7���� 9KO���z��
	������Y�8G�$��z���U��Z28�g�\�n�����2��ل':e.w�\��\Mˬ�� VVUb"F�Z�dvaA�2k}ZD�����+���x�����k��~�n/>KGB/p�A��k�,�T� ���=Y�?�����E~𶓙?�V1�@<7GC#}�l�d�l�W8�fcF�r[4�Cu��T�/��,�w����5��V�j�A���o�5�N3m+���6�88����w�"*|5�!�
E��S�GEW�BDW��	�
�)
�зw�W��:r�6�����7p�^
+ce��-�j���%�����|k�4��Q�������E�9h�y(���H�KWLZ�� �J�t{�u�ZZ/�ikGm�ﳖ7�b��e����<��BT��_6�������ѣ�����X�����J�`u)�M2�,uN첔�g�7EM�?O�l{����`
��K��������MM3��w���eּp���5���'������JށX�l@H��w���M��u�[�t���*:sW���P��I~G��`T�:�a^�GV��+��Wh���!��q�����ha��^W���j�Iظ�����B�S��K!dw}�c�$ �y�S#�T��� �'���m��6��M0�)W�~�������/������¬A]!r�x9 ��<:U������'�� w���W�~�샜�Q�ՕA9��.ȅ���x����h[8!8w����܂4�x�����;����.�q'@pw��wνc�?�~��z�)�jת%��
&28�c��1[	 ����`)����ȗlUk��e�~Am���mW��n��O�6�m�M�9��M]����]��u$�mH{u�h�Lo���	A��4�(Ol��9愼�`�l��+zI�Mm+�Eu4.�䯅��x

��5��]	��lq�%�� ym��?�:E�U��WV],P��C.:Pp�tI����[�֍�W�r���� .�GJ�OB��[p>�Ɂ��wx�	y�P�%����Լo�$���H�vO�!��Ζ�q��w����]���61�>�M^���6=yU��v�|��ٿ�$��d;_���%(����Z�4b�PN�q����<��Kc�c`���������B�	c�����^���-'�b>���khh�B��}I�����.��^��O��9�9~�=ٽ��a��2q�il}�W���Q>�#+�l Q�zh4V0k�~�����THH����h����m��Y�	�H���A2���U7���%n&�\�E��rR��`�;晈ƨ���HJ���J I��V��Q��"�7¹���'n���)x������t?���H65���؉���7̱"ꌧ���^��H�\��Ԣp����3:&�Z�q��N��9p�u~�Q�8�z�uP�]��(Q�\B�{~^q�e�Ss��Rݾ���- ���4hv��%^�0 ́������i�����ȞSdL�:n����K��~�r�X �]f��a���+���Q��$`f�&�i�i�>+���ޮ��>���y�%�_���X�!@����v�'^�8H
RB?)G�w�V��N�]@@�m�:\���K�k65�!�p���#MD!U�AW��ne"��-�2�mE��8O��8mA�Ot��3aic�z���X����o�O��5���2��B�i@H\���[S�vg��?W%M�-���t�<�GB���m�������R�p�p�iW�,vܝǡ����}Pg�?�M]���kW5�8�8�.'�Z� >٥���"(�)ƅ����<5�I@�Z��a|v�:��Y��-$Ε��r�̀v�kV!��.x��X�i�`���J��C��~�@�A6y��Utc�>x��r��Ș��!�"p�r��|M`���9}������i^��%�;��!w�|]�&��튀4�f1a�E����]�+ā�+=6˱ )�
׈�<V�۩�1�j�ώ��U����?_��Y�"�TB���1�;�ѫ��k+���U��TR��'Xa}`�j�T!ă�MvuV��t�s��Zky��6}]k���sˆ��Y'�u�Y�v�\��}[[^F&Ш��`�8�,#�&��������z+kԇ�c�d�-b��侞Op�g��$ݫ�_�}���,#�=�V��-A�������EݑXe4��#��CT�ȏ]��V�����k�_��j;;{g�U
�0+��y07X\���J�Z���Y��kd	�株<�+1Q��������9��B
(�(��(���a���V��V��?zaj���Ri��E�b�s�l�o[�;�N�￩o�@DNAàт�r�s^��d���V�f�������F����Ē#���̡��)��#]�4��x��
��1)���e!^�,�����s �١��Q�L�2*j�L?HSz1X������3Ho�+5U^�QX�V��riHXM���:�Q���Y��7�1,�4����c�}�k؄~`c�T�׍���t��[��{�S!�TW��ǄJ�oD��s!��O����d�%�bM
k�Xzq駛}E��v`�s��+�7��B������iN\�n��'4�Vg,�9����%KV@�0�
Y��ղ�_\<<��5G����b����y[ZZ����k��'�����ߦ�����ƫ��o�F�B�k/�;����Q�C@k����Pk?���d͉��A�D���eN�͛m�ŕ�`�����ޣ]ȉR�v-�Gu�G���%K��PM�y_*)<�X�f��Oe�|�L-�$�;;~L��&��Z[�:C!n���C��".�+�N^���-=��vC�L�ܝ  v���HTF�	R4w
���Z~D�ʼ�6��){�*i�|��L>*�~"�Jc)&F��Q90;�C��2{?��p����6�.B�sQB#9��&y��sE�����Yǝ���hk�P�����*�dfN�aP�ʣ,:.l^�;,͘ �G�K�x(v!^3�TӾv��=�_O�kW�:�]ȟEE%exZLVhu�|�:��XhmK����.Dq�U�sҧ��
�W@��~/M8�*����}?O0K�NR(gȁX���5���S�I���tӆ%v��<h䷙���ݻoˠǬz�mJRn_�o�Tڎ{�"��k�D��������:ffb����!�R����^�f�p��W��Y�C�gDE��[Y݋���め�O�@�k����@	$�?�z�F��2BvV���i@�l�<rY���g&�z���&�m��Vk����������oj$w�������,8�s��K}w<k9����_*]j��7�i�[�e�~���vr ��jL.S�-{���~Ű���������5RFKVm��ƪL.��7�9� V�
R*�3��������,�'"�/ˀs�&���V$�S�����Z��N;�X����˱&�������.�#����Y����)���'ZS�S�H�r��UDg�M~l�:�z[ [��ȉ������!��ξs���$�4P^��nR�{����6\�ϝ��R�>�}>����r�0+�Z1�8��e�û�p��l�s�UY�"�Oӗ� 3D,�D�, ������QXb�=�9t���چ������.We���4ˑ&iAˀ9^g��<��ʏ�]������	N�����5��C�5�be�k������Q�$E0j�_<Ξ���֟�\�jU�j�+���G˖x����j	[�ľ�(��ϊ�6c�� �iWy�>wS(�h��D��/K����
dĦO�]�yf�Y�Y���I�?��Q挱���腠&���|�(�e���%c�,1����� r�<K���L�̜y�N�{J\6���ԥky3��4�9����O���'��%������d�A8�s%�?A}r��*ܻ&�2g9O[Y�"�R5g:U�VJj�m��$�L󍫥�G�iTK�
��"�*�M�C�R`�g1��AF����� A�d�|���@�v����nD��*��n��`�s��;�ɶ\�C6�����ϼx*E�&�>egT����߈�}]��<#���l5��HEk�!1gm=_�׀�� ��Z��P��1�����tv��x�L�w�?#4�(��d$�~-b]u�aT
��c��T,YDu%�Q�돂�s
4���+"��Ȕ�6���L5�W���y���]�ݟP����v��$d����I?�����n�l�ݶt�J�u�����l�Ƭ����w��F��e�r���8�p�[��-G<��h9�x �,���i��Q۱�j�o�s<9�ƴ5��p{s=xT<�묁3Y��m0�rg�rw7*�#v1�G���1Vs�6~�[3��w1����O�?	!��a%�4�S���V��a���B�vY��B��s|�T���"*5�eg���A�j� #�ޅ�F@jІ�K] &>'g��ɣmz۾R��q����jXm���ۥ�������s�x$��u)�/3�ȿ�j7^���t���)U&��׬m\�j���|
�+AN<�d3���A%��.Z1���)!Qf�h�$[\{���$K2P�"[�QQ���D�tA�F��vN	z��{���~S�Ūn�Z� ��g+m��׈�"��k|�[`�Y��̅��;�gg���ՌV�TpѤYe�WkzYLLLi�-��##�7�^���(�2>!x�t5u��}�NEl��*v!��J=5�g2�ڔr����O@��;��>���2�]�ȋ�^�C��gʴc�ƣ���������Kp�,	�gu@�t>.���?1.����B�*i�/܃$�39�o�1>��gP���x�����&3l!�u� ۊq�2�؅T�dxp��w��K�Q��."/ב��A���~����X=hgM̲�\�2h~�0zQZ�]���z��# �+Sxbh!�I�OC
���+� ����w�������ۙ_�i72���3�7)1��Fh�b��iqT\:���e:����&��������)R�aR���0�=���u�<�T,�FG�L��3��Q��מO4;G������t*���^v��Ď�gÝ����R&Y&t�"]{* }�m�����E�����b)h�Z#54�̙��]��y�������¾���6;��zf��-�4k`��z]�J�C܀1e$�{#㈹z�2��`����X�eo����>�,�����c����6���\"��jk�,�=�����uH��@�����}��y���Qe����>��1+".����Ig~�5&Z�uDڼ���Cg� ���X��5+�v#�X	T ��ԗ�Vyy���p��APf	y�  ]�lΫ������ݏ��umw�Tj�����Q��P26���H�Ԕ�S��e�~��O��яfK�÷c����h�@WA���x'ABE�8ȡ��w��@0�<����0]
�꒟/6���$F���7?����g�M�  i�d0r��h4\�kҿ KJ�^x"���2������ld��4����J��/�%����	j��~)�r>�)$o�l���Y6���*?1]Z�y3��>b�+d��}��A�����`]�����{��/���%�]$������)����ɢ��
�(,Pj�WB��7���XuxZړs���:L���Aq@y�*�����,ʬM O쏉(f=ZB��Ꞗ�yzϓ��G���r����D
���u�~�P�Z	M%B�Ne�Z�}�`��?��:?Ϛ	V��츮�Vw��֜01�OM*G��==m�,V�BPI�d��ź�y_D��͝<v��<��^���?-	~���;B��yݶKe�D�`��ƬI�@?��ґ�G���,���bDZ;b���[��<+�K�'8o�{1��ݗ�U�'��w01�{;���x8k9��1�K���Pe�D�zkm��\ܚ/S���_����a�e=�S�$^\�N�mPJ���C�y��x�!C�\�n�p�C��9����\�R�?��0p/ى^�tpQ.d��{��񢸻���Z9Z�Q�kh���3[�?<��B��W����vu]c�y��/Ӷ,I�����a����،WL�ۆ>��{����
$Yu����I^3�4�G�Ѭ�Rn?�Hi�GG_��L��p��l�;��3dpH���Nߝ�e>Ү�G�Inl-�V��c�	q	))�=ϖqD���܈���J�b���C5�������r a��΂���G����l�C�m1�u�E���q΄��J��2bc����j��.@���ZcZ�ș3y�p�t����_��2�<�S�zsSS@�ȷ M]<����2���?W�"'g����1d?Q/ ��Γ5����K?��I��%py�0��r��3IG�{����)]hHW�a96v�h����HVHIHfѰ��Wems�D�*���٦.U�����݈��}�l�^V@#&�Z������S,S�K��-�6�f_��|�7P�X�M�x-`!]�C�c��λ�1���pū��PE��N�!���R��$���I?��K�E�0b�g\{:<.����������r&|۲q��2��) Ή����GI��t�*SA��	�Ǚ�VyʉV{q�3�V���/�6�P֥�B����C��`ҳP��^��,��:v0��q���	�� D�Z|�K�!�<�X�b�u��:�V��ۈ�#��a�b�j��Q�x�	��Y�,W>��*=�`Ojhb�������f2�w�xfabј�.APEY�re�L��S|dd[6>/��L	#�&�+��p�����k

��U#"�v6v{����y��2QѲ�1��yg�aJ]��*m%+��WuJQ+��D�!D"�P0�d�\ϝ7[r2����(�b;9y��
.I*ɲ`��0pC�%��������m埭p�s�mPy[�������՚�>�~Ĺ��YȠ�trM5C����T�ﾩww㓹#�:c������aYM���l��Yд3�k�c��u�'G�����=�CN}(�Vx$<K+V�TZn��*�pA6ڐ�~'����e�tN�1)|tF̭d������cM�_���1^E̼��p�xU���n;*����n�+���\�&���9G����"�S����	��5'��=9�{(k>c��<ݞ�{{gF�d+-�z-��|/���˟fSGb�(����?��={t^F�u��d�$��$�Y��V�#���I��($��M(wv����S6f�$0ȵ�rz�?&<0�^��>���G[��m����6��Hn����kb/YsX�>տ��j{����ޑHc$� h���ҙ�t�26��k����T��\�,;�rهk�?��d�*  ��2�����/�Z�d�<��"��8^��eʮ���
]a�XD��?��H���N��d��P�Ffg֤����Cш�/6\�o$���uQK ��,��BBoTq�����2~�t��!��K�,����{�@d���~Hh����~؋�\A��}�@�%}�y���^��;\��V%X}����@��xp�,� ���"�(\ӻ��ia�>j��e�d�j�x���y�d�hX7�y_T/�?/t�U��`Ws���
�������o��7��jdd��᧍��{@ǯJ�s
����v�}i��c�+�v�<V��Zyyy1�i���P�"�渘Sn�X߶�۶�.�����򊊱���YLI�0��+`�u1Y\Z��8x��w���E���XD�߸��J�*�0	�i��o?*�S��Wl�eĔ��)���c�=��ɖ��I�>�����y�dƒ�sO���{,���ր,h��6�gk�|Y=5�����F8c�Qfa�ͩ���V΄h�B�F��b����}ߵ�$,���h����h$G�����mD��
>u㣗lO�(K�7C�%~����{���i�D����_B�����|8ƁT�Xwd�7+�ws{Ol�ﬞ�s���x�G�Y�:�x�)��������G�Ld��@�����?��d�w���
oµ����%;ML"�\�-��m�H���r�~�c�XPr�h��WEf��߰�=��o[�ۭ��Rz�?U(��yީ�U���Ŀ�lמ���nh���.	�Lq�qd�12*fζ��֋����F��s��a�7cq��'����[d��f�eU��IO�?�����9��DZ��X"���ReIC�$�%��?[Th �l}�BNAΔ7̯cC�wcaZ���&lD꾽,�=I��Ԩ��&��j�l�5�T��;E��V��}1��F�4�D�F��Q��̯ʽO��U��L��J��3��i�%���[C��0	ҿ7kK�����*L�X�wt�8_�J��z��E	K:Z�P���Q�͘dMC���GD�o����d�EA������ o{����h�a[���U;F�������NU�K(�G����63�m�����%�/)#����۽�K��i�]�\ 9q��'�@I�"���o���-C\	�����0D��R�\y�鳻��XŎ�ʲw�w7B�ࢇ��p�y�&4B��!i�5)[q3�~Gb?�"�+��e�<�.�T��/0r�.z��
ꥴ���[��{�P�7�^�>�����j�I�����"ݿ���k����FO�^�2X'��.� *,�r�/��wW���:�����YU�h�Bo�όhr�ޖ��H[j�֯�&��F��}������F`�}5�~�э|. kF�<��''��=>@�^�����Xs=�_�|������cv�;��סcYC�eկջ�#�+i���YUՔy��S�@��4�l�S������'�A�J��i��<���l)`;�;!$�����&�o���$ Z�j �B9�9G�M븬S�؊C�~�&��H�ùM�<m�����"��3��;�1|0L
ww""Tԋ�p�7zF�V�)�&gF*ǐ���r/��JW�.�u5�8��]�@6c/��e��0B��`d��=N�#�9�!����4`}���P�Fn9 �F#�J��w����r��dƠX�c�7j��ù�@�Nl>!&y>��C�~��C��L��Mn����Ky=�յ��×^q���N��L�.A����8G��w���Ѫ6d� j�x��D��ف߯��MAC�1-;��|���i�6���Ձ�
]���(���w�G�����-g�wR���F��q����J��b�W��9�[6��I��ko��%�fQ����-�NKK��c:*sN���2��0Z���%6�e*��w¥���Qp�'z	��睧�WNWȟc�`�Tî�'v�A��i!BX{ڑ��F�m*8L��U9|}��ljO`�����L=��
d(�4~��ŀǆ�z������)�ı8Es��Gp���1�([D���f�{��װy�V���("��^&<vC0� [����̥ ��NA��e��������ZV*k���o/tm�I�6����}N���ݦ��������#��[(��+����7�8�)�hQǨ�%iik�@{� Ӳ��mQ4f��A��kBH�ps��φ�������Kx���f+��$8,�pE�[�P����ZϙuTK�7�����=�f{o;��͑D�������J�=_�_�3�	w�TMe�J��[�e����ѡ������!���{���$܈3�����=w���~��� �o(A8�ح{I�ѩ(�2�,��=�
b����с:�	w&ɂ���a����RL9L��@�3yK�J�|p������Rq��^��~Q�âa6�n3�p���y6v��y�imc���cQ������Wq��c[h:��<����ݘ��Թ����Sm�]E��T�kס��Gɲ{�ٙ�e�f}�¾��ĭ��o����1}8 
�[����u��w���v�u�)��4ye���s�m.��_�������U���Y��$�-�qz��Ļ��p͑������:~u���c/��~l5#�q/��P�W ����uX��� ��������������eŭ�PBv��D�d�����cX��k�*����2�t�����{lH{\Dܔ���"�3q���E�O(,�_鲊�Z3;�7�_NR��U�^���k� e��|;-Dh� �f�f���/��^��
m��u��:��	S(���z"�d�j��z{=��^ A��0s��sF���I��gj9f�������(N�'�ƹܵ�g�O�Ј��Yk�ʭCUUk?�wκ>cU��H����߹�������߾������c�)=�9����>x�q����V��d�)��������~[�}>�f�����>W������t�M`�d�/:�W�
�bW�R2PL.*�&J1ĳh�J�7��]Z��R��G�B}�9����׌;Ԓ����S1�p���1VO�Am�����̊ވ!Ƈ�hl\�lRKi� _s�z;1�H�L(��P�d�4�d3�R��䟨#�3�Q5Dk�K��#i��󴤇ͳb�FE �R���M����PC���c(�sc�
���,}�X<_��lN3��� t�^�>�e����8h�n�������~�eVU���ş��88��_N��u;��1����4JV��UQ�R�Xc�qq�`Ԩ@�@�A0Xk3�)<�Y#_��}�i��#J��"�������8��U0� [ܹ�&ޖ��'#��f��ī�� �^���A�)��rN��v�w>o�{�3�6�_-)d~a��e��&_���iV�cT+A.˹O)<.���n������y�������A7���^��-���
�J0Z����H0q�cM�\���פ��`[��#�0x`=�E^>����_q׿��@;����j1`�	%��(�S/��/�w�-�Z/�O�ޗ�?g���(	q��NS$ӿ��F5��P"mk�K֗�1�Ez�;}�Ԙ4��u�@hJ�"cB4��<e�<�PD1�jb��[�T��isk�`8T�h��-}#���;�����c��cTa�wA{��(�sv�;�u�I��5�Rg�?X��F��9�P�WN��
b�����y�H|���/J���Fд�Ķ3X��s��g���s#*������W���	�ν��:���#���00�Yp��8��u�ys�(C~�~�8�9�*w�:����9����g�_������Ŏ�Ɩ���)fx�Q-�|Z�~X�*<���V�j���4�/�X�B�0�z��Y�����U�e�u��Z���,"aQ��?�`������h��v�<��j��Kn����S�;ڪ#��	;C;�+��ǫ�s84��wi�(O��Y8`�Ȗ�8�S����oó<xJ6����e;D�깞�8s��_r��=�$g&�Ӣa.�����nL�0K~W!����%���@,�x�h4��f/�<�ʼKX&)����f+S'I�lI�1W6D�����O��3��S\����r�Kn�݅/m��E�.����ӄY��P�
S��^�k�����u����B�<5�m�L�=&��m�s�Q�>�%�!��cXȢ,K!)���'�b����c����ޞ$F �LX��e\�>^���剝O��9I��<��k�ҧ_t�j9����9�����_̓;��S�ϖ�W���ze�<�z@($��i�ރ_�y�܄�A�{�$�Q�(g罄:��)�T0b�{	d_��Qxz�`9�����I����Q��3��$B^�������r��S�e=|
?�l�K����YTJ	:���>E�Y��L֌�Z�Z�	7��6�WϞ�ș2^�jэ6+��&�މ�B�1��|�%�k�?�8m������p%��b����x�KW�?�G�o,)��C�_8aK�sp�l�!>jC<.]�\����ٖE�9/��<���>���J����h����&N_N�h����Y7k��{ަ[�CoAX���4����4����}F6#gϧ]�s��i���$ą��b[d�������^�6����č+İΣT�U}�� 　�r,l�� �+�Jk�AB¡�z���68��J�G��,����*���_�2q���gQ9�2_��cc���:YZ���V����IV����	j	&uڝ�7UW̾qA-�)�5���2�'Q��.�><�*�!���Ybw�`���He�
�aR�D�E3.�m�+��۔E�e��������Ыnq����U��3�Ie��I��La�O�m�e��iJW�-%��_&c	3w�{�;���-�+��r��D��բ)��Zq�Xg����Y�E�l0"FQ��	Q(�qM�t�4l���A����o�������P��y��J�'Q4� ���)R'-��|�Zp���%�c�O��/m�tjWr�s�S7	Dd�,�����:�\��&��$�v�!Y�4���g&�yIs��u��Kl�e1��tC�y6��R�Eܸv�9��ع���k��ǈB��me����::DU�0�3f��]�T�0�V���aI�t}���f�p��,B���voc~�@F��3@Tt�����U�@8��
��pu��U+=W����f�&�����>�����g1�L��1�1b�틻��/�7��%J���Q�J�4i[�*�\�y��WaJ/����ǀeH�~W���G,9cJ��FO�0���H������/��Ru��W{�NX
����s�z�L�Èѣ�Q����@�h
��4���RD-���|*.N�%(����=�6��Z�gsQ��Kԋ�~�'N�� L0޴���;X!$���jW���h�~g�m�e��/ <�;?D�Ͻ���;l�!��*˷�l;�R1�!IZI�4�4Y#�5Ő��o�Y(K��[a���R|���F�Se������;���}.z��X��5X3�S�~�\�:u���"E�Ȟc"$�=Z��	7�k����_��7G��=��m^�\2���T������ܩ�9s`.�����6m�I�]�萁q�L�E���/F@�B�Kvxt��U�Xy��l�	n�i~������U���.L�XN�a���F=�-ܡ�����A<"��5[��m�`Ʉ:�: ?���iy\��]�_���L���{c:4���Up�\��;A�<sP�t�#�u�ߪ���R�!%�&�
��}�#z����%�wV/K5����Lq|?���
������Ӂ2k�)�
~!��L (wq�#�Sn(
z�m�a�~�=�Ccn�-1�o��ZCK4�ab㡣������Ȟ��Ǹ��� ]�J����O�4c��L�\�<��{7������h�ԃ�U��;\y(n���_�����V��a�TbE0ɪZ�"�&?����ό�[���=��>�Q�:�10�*���S�S���΢C��!W�Lʁ��\Z�c8���S����E:k|z��i��oz����eݴ��80|������mV>�Y3|��Ka\ ��6"���cK2�m��w'}O����b�t$�����*d����tX�#�C�醖��=AW��Lj	�|�
BO-����]��Գ:�f�0v��E�8SSz�㽒��tj���Ǘ]�#J�_�k��6���cP���}�=��2�����������pX�LE��iu䬋Xz?�xʔ(LW��1�:�t�}�N�᎙�˪U,�`jX��P΁ŠA�3bF�"�:h�L�)����[<�uk�<W�x��1iU����UT��f�^��A�v�F= X��b��W�`o���bA���!�Vs���;�b�k��;�m��e�J�yJ�j3e�y�kԞ+�ς�)P��Cхd(�u!��	��"��]�^e�{���+����T��%�*��g�`X��C�W?�3~��s�lU�tz�B��Q2w��r���w󓁀�-Èw������K�X��L���M���+��y6���	|���Y(^"��]oH�󽄲���G�2+X�?f�!T�|�|���<�s�g]!�F�S�����%�	��[ܾ�3QT���U1�H,Y����`;Qм���IsW��	���j�o�H��F��O����MJ |�+r7��~���������a7b��K9��}�"��c��)v��rO5�i
D�j"���.J� �����ih�����0�=˖��=�x�kh�-�̲9��ofo�����y�4��1A�m�����y%��L	]�������#�>�"�΄aҳ��	G��J|�7tI=�yl��U;�X�;��>��n�x�vѾ+�E�`�>
7�5WV�*���sS��`۬*l��% ��q�j'2��,Ӭ���h�hX�9/�2Q+�O���	
���wS��A�-CҰ�;LP,���	
�x�Z��=�������n�{���2�>�� {>��I�yR��!�v��[�Z�{ާ@�]'��nL)�#�D�dxik/��~��Y	����C�~�oh�K�
��1�������vd���1�R-
�=��k����.[AxOV��>6����QN��)ji.�p�u| L�K(������*�Z<dr�Hޙ;��'*̢���0�b^� ��C~-�O}e�<.%R�VF�z�y��ËӀ���ğT��0�#���33@=�>H�'���(mV-畨֐KD�+9�+���oؑ�w�g��������'�������M�Us������|�h`�dEB�Q�V�j����9���r�3u���f����^s��l�?��GH�zR���gQ���3��2s��|M�g^�M�@�-}-uH�(ѬBB�*%������ic��]�g�kO�~~�w�h�P2����/G]��y��1>Sn�� ��$��,i[{s8ڴ-�tG�`7�	��������>��	;ղ�3f�ѨrI�A肚d�Qh$�ݔ�bc�2b�*�I{�k�$�N��BO��)9 ?�v��P��0&������WDR��Dn$��M'i+��hȞ�KD����hl��dC4wQV�]���1[ �b�A�4i�5o>Y)�O�ן7:����<%��c��UH�WB��錑��=��w�,�5c��o���v�h����m�n+��2� ��U+�͟���9�[7Y�}�gf�@�N����V����+�jmck���4x��9,�f68����v������f��C��QQ� �|V�^jLoF0�Z>��	U��J���f�L�P��1W�|��ϑd���������a	E9�lG���!���b�--���#6�sR��UY]ë�a�E�%�?&C�Q����P&jߦ<�Q��+N
\�zam~D�������'��Q{��F�4���v]�kn��e��7�K��JF�����f�����;��^[��q�ly�##�$�s��s/�4�{�:�GY��=��Qͮэ׵�҅�E--����s$�G^W{��/�R��RA�g�jd�P��]E_���9
%�����R:>w>W؁�.�w(a�tu�m]qӖ����.Q|���:Ós�Z���Y�>�����FX�N0���d�q(�}Yd7���<!���=�0
�&=���I�؋�3�e�{�s)��WO�80lQ8X`ɂ�=3t'f�'�Aݕ1��ۃN�Dq��\7�����I<<%�<������ׂ���U�i9ā��e)V��k[���S½�:NU0��%w�"����N��^^�|�V���&<w���$�g,�J!G&lx�R�x�fe���tT�	l�������J��t<8�L���6+r���ɣ�㒁R ���z�lP��-����V�B�\qu���<n�b���7��TB��Ѫ�Ѻ)��r��߄�z_�&�>��.�N|�!��P��߲B�N0�
�~���{�\�҉jwY���O�eM�%x�'���A�.�IV>�̓�	�+��#��-� �!?�,+'�(y6)2}y��� C�Y�z�o���=F��9�x�g�t����n�.���mD#��w$$�{/%��LT�~"�G����x��o��.������F�d�������
J"�&��b�H64&S��\	��������f5rEĂ�핀!+����w���GЊ�[!�驤i��tXa�έ
��%�Y��g�i���9�2�М���qߍ
n{��ߌst��Lݭ5���+�U��!2,@q$�	�q��o�$;v���s.�t6p6�q5﨏���Y�}��)ݮ&�Q*��F�(w�7E�ba�5ߘ�P�2����A،In��8���U8w܌��GҶ��}����L�aN�����$�98Ϸ r梜(�n�!����p�vV1��ޫ)`�)�N�d�_{1o��l����x�ZY6N��^7%�	���s�y�t�3�����Z�|�~*6�o���L�u؟�,жS֢7�����B��T�gcR��!�j/+t,�Vk��Q�OF���x�`PCW��0��'Ö�3��PQ"�b�� ��f"���I݊����{vv6I����#�GRT��l��H	�"�2��y�dy_ }Z?v��7`e������(R�b�$X.�e��0�D�ROؖ��7Ȩ{dJ�.�6�gyꁌ�k����@����e4��|�ݒD��ٝϋ]y����j�E�,�Oӧ��)co�H����:���22�O{�+nSfi��6��?�/�=?3�����u�����nS�iD�����&r��F%=>3��6H�Ӧ�u��5��"�=.�b�+	ל'C���_Y�G�]xp�#�x]��b)\ �Ie��ژ�;�)�7�&�2�В9�_�Nl�E�.��E��e�H�9d,I���Nk�iTm���&����y���EO�b�'vߍP�#�3agOH}B�W��I��c�o��<��I?��s+Y$�k´JXߣr�g�xH��uI�l�����G�y�TG��?A��81�+�� t���{�s�p�!q��ۚ_���6D!�������K�h�z>�����x|��ȴ�{t��Di�!�����S��`���=��3L,Of\1�^�i.:�T�*$>��IԺ��;���E�A�2222�4t�t�
)��x�l�b�ڟ��/�Wa�����:V���\/��N�-08��������Qq5M�������dp���Np����������ߺ�ί��Y��wծڧ{�zF�L�N��r���L��̘$���)�:Ԩ�v��7���8�z�6u�V*A��Ee;5bHIu�E �p�h��%!w*����N��T����}V�[5�?xO>^k�^��Iܒ��i�.�ݷ�C������"��w=�P+R��}�`#i:�z��w	ɦ޹����Y���ʹ-F|X!��'�0�哾�-�i���C�6�d��2n�	���J*�X^��!z0����BT~�ʒ���X93W��b'A�j9�u����t}	�{|.]�~d�$~�X�
�� Wu��T��n�FDD���=��o2,�^=5;kd(�x�7loG4�RAnɤ=1Gu\����#$$y��pǌ��v�������}|~�W�c�@��3�o�m4����)%�˯I0G����b7�F��"�������P6�T���/9�~:�0�@�ÜolQ�xZM�	�kewH�ީ"����L�@j(,O7�f�y��b��y@�;vt�ެI<��9M��j���X�������UMU�۱�ko g<�^��Ŀ7S�.`��s��pNF���΀ N��ymvNN���z�D3���802�kaq�D�fY�vSj����(��z�-�2�rFS��Ύ��q?�S,e�W��8r���7�篓ȷnYyj�WGC׌x���v�*�n �A�������ظ1�ۖ�aF$�0/��;h$���sj��4��N���y-Dk��-j��й��\���~m3[#P��@���J�jX��'ߞ g���-XAc����˵� ;��Tp	�3���a{a�g��I�|�{6�.�3�:��������XB[�B	��Y���%-��Aө��9/��7�r��#���^8��Q���"hk�M\�P���@9�:�85�(��|�2P0!�Ӆ`l�5>	���CT0Nq]C�&T�W�~cȾ���Ƴ���E����c��s�{~T�sNVz/G�5�F`����콓��+"� B��c8"�'�X�7@7{jji����0�j���OҊȭ3!��xŇq��H�Za�P�~c�>L?%ʌ�E�>�TX x*"��/f��b�n�LN��<��5K��g~-�I+��7�?�{�yM����y���\j��Z ���S��%0���}t?�+}��F8���3 \/Q-�,����i��J���L5�������T�]�'��XO�a��f3�y�vX��[J��!�in
%�Q��l��Uc6N\��(]T8�,��V���q�>�␬�*���ۅZ�X�`/gHs������7��7VAE�a��'��<���ӗ�p�4 �@n��c�	%�[n�Jxlj{��߀A~x�|Q��Chhy�E*������6�k��d�s�"�|�����1�:B�������c��W���i�"��d0hרn�w�΢ߚG��ֻ苗��iB.'��.'�I��»���4�Ͳ|�Z������#���-|mCj���HHHU�B��#1I�E7~���&M�r.�vR
�t	PP`�W0}�/u�HJ���KP����}��t�-�l�_���)OI�r6,��y��mU
�x���n��>������,�/�*kZ�;�L=Ζ�wfҦ]V>iQ^���Z�T��~vMJI�0P�A��Zs}��]vZ�?�*�MS@�(���$@	$=�>^��	}�)fH��&�{}���N?�C�&<�������_e�i�3����K;��So���7���ab����c#yE��*;4�\';��;>ׇ�5�٨��wL$�Mkj"a�&@� Zl$"!�����l�4�+��My��L�j�.Ѣ��j���E���m���i��qF��4*�T��6 m19 �]��6۟]L�y�yO{�*x�z�,r�(�X^�y���o��?����ݼ�[�E^r4v������k���W��>w�/]�`�rN������B����we��� �}@������$�"iLjUz	�`!z��s� �/Ȍ����J�2�
�əaa`�4@S�\V�|Y?�@���G}�����7�9僲���j��6l�[Ԡ-�q{\l{���e�K\���f�B�`#Z��<�`��U��w��]~�wp��Yb�\�lK�s!C��?�En1�[��G'ځ�7��_�q@誐���J��-x�P26EB "+ x�<C-p���3��R��]�|�,%P�q�<.
+
Y>rǹ`Tݮob�C�9K��#;F �#��0��c=�<~��-`is�Or�̪:���(������|����ֽ�B��<�����by�B�&���_�-���	��*��(РL�_(�(�,s�de� 6�l&ܷn�n��9��x����b6�-��7��&L}{?hP~Y?OI����Fo�'Y<��S*�x����2c���/���oΞ��A��WG̢���^qҎ��������qg��x���偕��ã}`�
)�<r���4!���[X��;kg��yFǶE�}P1e{�Jw^Ǜ��,64
,A@'��n�4�d�BW�3�,!GU78ĕ/n�?��7���g\mǩkh(�\i�ti!J�Nk�j�w�ݬ*�!ن���q�K��+D3�p��:Mi���,�S��[�Z����"2:)"�p0>&���1���C#"��d˸���dD�":~>y�HC
 �
�df��
*��/�n��4���MFh��F�u�
]GUY��h�#!n�9u� �{RZ$�	����)�,}�����(���};,#�'�[��q�����t�i]`�^g���y�i�
�J�T(��wYh�^�n+T�3S�����Y���S�nJ�a�
���c�\lC����7'�o������Z�֔7xY��~�L*�{��萜w�	��o�.�׾�y�, v�P�=̿?��ݾ$*�)�l�Q�����԰:��1�?1�1B��'� X��h���l���C����7#g�+���h&�C�@�J� ���U��4N���JU.�6!&.�?�>Uڟ9O�K]+q-_�����k/z��\������mк�F�Y��r�F�w����)�阢��o~3��n��n�~�����M+�v/�P�\��,��������U}��4��Sbo8��c�-����I�혭M����B �}7���/ק�]WR�?V��ƥ�ڞ�hy�7c���[Ճ�����I�>����/-��!�\���kkk�d����Lb��y:ވ���v:GȦ.9�Ւ$���zP"����j?�Dh#
��YYD��mL��Z�C9	�my���L�+��3���4��6c}o�T+�d���v�2��^u��~G�i�܉�K���$���ښ��w��k�˳��/�p4>>/>����X�Zʍ�([K8�
��NM�&!+Ҫf�ks[��o�U�1䰎������p�,2��K�8�:������z����X! )���?���yĢV�������i�V"{�c��^���1D�������]^�+׷��(�R	��y��Aڎ��7�(�����|\�1�l��jZ#V�r"��)��/G��̿��M�f�����ئ�4Z���;:�}gW�T��n�U����%I�tfb_����3�5�[3������X$<�%"ަBs_X��T钾1�O��}cH���;�gl<!q�6��/B�c��~���8E�$ד	
.��W�� 7oX�fi(?��i�1��O:�&a�0���u1��$����Y|������.��.�t+D��py�bY?��1//���b���x��� T�!^/+�_[hI0(�T?�X�Ga]��\��R�]Ż�?^�{�z�)hk{���=L�	/*R�fdh��D:v�ڝ��M�Ԋ3��J\��g�Ĕ��:�x~����C�0u�0Y����4��r��&O\n����@��|����L@<��K���!3�u%���}�)�9:����"xN�)(\��$��t�Q���f>+�rK�_|�"`_�����Hk\�P�fZ�]0��{A+��-,g�n������ucup��D�>���q�(CjB���t]��7"���+�D����}��a�l'M^�?�ulT�.�{�
�}�<�.���҆{�amȞ1�	�+)uG�D"ܿv�#$%��e	��~�0ԋu�x�ǂN;�+$ŗщl�dM�����t�B�j�=-ahh��-V]ͩ��=�L�!@:_���4q3�(�����2gX��Z݄�e��E��+���(�z�bX7��s�+�畢��U��F�Ҳ<шW`��y���J9�4�\�����ox�(�vH{A��JH�W)O����ݢv;0F@�������:��O�mP�������=���P`�9��r�9���5@�W�G�	�j�um���9�MR�J�}L�~���+V3���w�Y�J4[�:�+M���=��j-w�6�Y��?�g�	�n�NUW����W�Y}z��@I<���������nc���}�MkF��4.S�D8;�ylt�+����;����3�f�̓�&�(8����i)�i�hŰ�~�?s2a�bW{�5���K����M2C����)~{�!׎��NW+f�T;ܮf�S�"d�c��s���Ka�Hq��������C�
=������
���Rk��d�l��G�)Y�����ħj�&�<�g[eF\���6G)��B%��%"~"�53�	�������Y�&�1�ɸi��ӺB�c��}X-�ʊ���Za��)A�V.�s�w>�b���,˅?���G�$,�>���s��܂
z�O���47R�j�5��􌼬�Ç�����C��x:o��cY����Rm�iY��4����T��haڄ�Hu@r	���\:M�ԙf>N�n��ܙu���߇\����g���(0��8$�l�Ē�CB
qNL�����4j3iX�!ŰE��N��$��.?��%�ᒫ'`e3�OW�\1��t�vn��ֆ栮���� �
�yڸ�Ğ+�Tb4�]a���R���VaD�P��$���T,� �N��_�-���ş�2N�Pݟ|��
����
�v`O1�E����e��O���&O]��u���b�zFF������3���/����u��]���뽸����;¬~'k!6�0
&c�ؒ�,[?#~=B�(�G`��M��F�4�t`��9\��A�{�u9�85��=b\'ʭ�I�Ov)U��Q��&K�J�u
��W;�r���1�޹׮�~��7���� �b��_���A���2$؃�ƍ�̅	c���p�7���!�Gf
�=�EF92 x�a6nQ6 L"�sV�Jn}��=�d�̽�I���V�l������+ WW�,_��[� �NA�����>ir��� ���s�u��r&����
q�?�,�N�w<�Ե׌�"�)uB-�6�efA3q&k�e�'ˬ~&��v*�.=�o��.�k7Ceu]MD&��dt�)d�_g�\��ku"pycp�g'�i&Cq��Ki���C!���c�i0G~΍��ILOu���Y�2Z�u�y[�	_/�e��P��p�C�X�!�����˪�r'�5C<e��l���r[�~�ڐ�:�����������P��=����.�����	����W����m�V=������;}a�����Ѥ��l��}��?mzOe�ʕ-�����ow+*�|-)�ʜ�-���L��5���5�:���4	���(ӆ�V!Y�����4���l��/<�I����4J[�:.";������к	���+l���R�&GƓ���YA�����y������R�x����~d�N�2/}8�~G���G�m�"C��!�8ٹA�12�3.��7��S���l߈�t�\��č>�u{���V�d���!��\�����r��÷�CFA�IG����!+���ei��D��Y_Ї��M+eu�)~h.2���"2���p�)�� ;O��g�w��5��������=��(��=7;D�Tr�<3��p��n��Wn����2��^Ly�5��*� '�Z�f�TƘ_�D�?Op�N��`��d:��ޓt�L|"Ȝ��(Q��k;o�V~�4xc
�f���|����\��Ġ�����т��Ɂ���> |��#_�k��D�����&�ƍ9���ɻ���l}g���k�čA��t@���ô�	ĜvK(d��M7�Y��}
E�I+�8j�Hݟ@��]����u�D�㏨R2#���f,z�*Bw�V�����⸹e�Rbժp�m�A��u�9g�$n�|����3*���g�(X�
�A9:~$`(��77'gMI0l�;k�X89�7u/kT(*��o?�-w��d�צ�WST�ޖ���oU�v"��"Q�l�cR޿$�絏=.�P��=a����Q����ߗj�s��m��p���ŋ�ms
��"KaѵB���9����~��íoNkX.�R6�LN΄����k�*�N��pܜ�$�x��|�D!�rĢ�s:�5x�Z��/�6�X
����eR�O�����͗#?X7L����/G�bT��0OO |Q���G|�=߿�9g�>�x�bK���]
�������!�߱��L��i2t#r5� 2���?�j"ȃ'��/mW1�pCz�|��d��0���LV\��l�VX{Zt��rno���'x*$�@��&^���)������jO���'l̺M"e��d�BB~gA��X�Mȉ�Y Q-��v��!�-O���Ӎ�-D3Rϛ��BZX�<Ib	��e���kL/�/�%��ߖ� �-J'�I@
M�Y��O�22;���]DcL�֕Mx�SIp����Z����<�q(
R�3�:��:�c%�.�,�I��6��!k@�-�Q�$S�+�j�d���Q��)��op�ڲ^ �S������h��I(T>��Έ�0]��ܨ�v��kj�^���}5���8��{���5�C�����Y��ە��څ���(Sl����욛�+�o#�L�:����~��x�F��xܮ��57f��~��}D����u�r��1�)�x�������}{�x��y������=����N�Q��7i��d�X�e��c�5ڿ���u�9P�deK7�3h��9�+��IZ�vC�	:���� cˬ1K��2�!�b���F;���j�-蚮N����LS���H�,�����㹻�9h|���x�i��q���bM�1 PD�9��צ=X�K3m,����|}���l!֎���!��i�J������TPb�.!G-a}é���� �1�z :p��"m�yi�X�$��ƭ��*d�RM�jҧ`1b5��ޯb�ء�\��1(���y!)�{Jt�+$R	.��-��mBkpƽM�ښ�1�6��;מRRR2�	@44..�6}�8�_g�WC�W�{0��hQ�,��ӿ�G�k�7�Bb�w��[_R%�P����ed
��n%�o�|~��"]s̃�W�.ՋkY��k%mcPM~!��sP���GH3�CDN�Z`C�߮�?+U��[�&���9k�������m�����`��,a��+^�լA%g	POəS�HI��CŐ�#�
# ��(L�/��.ɬM|#fL�v�G�2�E\LH�m�/�Q�!6Sc\����W�Ǯn��`���.|7�q�}�Ռ}���h�Z9���o�Bj&��~�H�ؒ��f���S:^���̈�b]������X�$1O��uݼ���`�iY�m\�|Y쐑����y��]���O�X���H�H��}�uX�NN�G��P~�,g�j�Ei��E���z��_u�-��A�q�eV�]�X��*$�g�!�,�Vko>��f���ڲfOU�Ū$��Ul�r(NTP�� ���U��fJ�=\u��7��aY�/�"Kn#�a&�b�;	r��c��#���&����t�����;�a����,�;�_��7._�G~{!�S�f,��TI��K�$V�v�Wc%�;�����0��n|�$�����
���_Rm����v����OS�,��ۚ��1���G?�/�;��=�Gd���S��}������^p��E�Э���N��r����l-Ѡ�UJW[ܿ�T��H'�s�i�X�I�ֵn��X{���t\Or.�7fKw�A$R����&�v�$ *f�Ҡ����_�o��m8���~1� �آ��6$i�7�I�TI�P�*͛�g��?pܗxۿ�;~��A�@95ܰ�ɳ����@N��P��0�;�f;�f'��Y�?�˗,�f�-lX��L©Yn����0E���8�4��Ya��k�^՘�]�j9�EYK3���������MQ�:h��iɫ<���ۉ�}	��-��k7(8�ӄ¶O@��Ɯk�Q2Ѹ��uv��X��x�) L���7h��7o2�|�_
Nh���E/�^�mo`(:<����uԓr�rxT]�w��eV���Ǣ�1)�y�"�"�*Hv!N���F��2��"(�fo�̌$��
(���#{�0�X�<�:�8��u��T����{Ȉ8�{�˰c�K���S��y'������8J'�y,O�e����hX6�.e������\pp���,�R��E�Hi�P�{BDdD9�<7��";�(
&�H'���?3%�%vǝ���A��G�e�;.Ν�@:���CM�/k� ʍK�����ȯ���`9nY�qF����>��K�b;�ZA13\A�Z�A�4L�S�m���dD�V�C+�Z���t��I/C������6:�J)�a�H�\h	�o���`����d�O'�8����Ao/�Sn_��(��=�O��:��^s���ֱ�ԍ{����}n���A�lc�^�RO7��- � ���qF����R��*����%�q��r�U�pE"y��
��y3����H*�	U_{<a1]�r�H�͚����m,&������@Ĥ���G�(��i̽שR��-[��S=hY��I��'F�/׫{�/jr�=�S3ѭWP�O4��@VҔ�˫a᝛puŽ	�u'�㠴�?�soT,/Nzɧ\	�a	�ߝ-��d��r��*��_8zB��L�7���za��z����~/slHTo�]���8&+.+���!�,L�~���</�ۭ��a>�}�x�����67$��.xKۅ�2ݸ��x�1��-h���ZH�ڤ�q1|����Թ�A�<@�1�?�ҥ%�j*$�����0���]��6P��p�J�`��o��./5�$Ul'�|9����FmxhpܜŜ�3�VmD�}�(@��q�S��C5�X���q��8�H�^�}먀�Ǻ?3��dx�ʽ�Z��~��)H�{�1c�σ1����>��Lghy�}����2���j�[h�f�])�>H���G}���>�CEW�Шb̠����`�j��w��� �\����}l�qq9���7h�;x���
��%���+G%��z�"�I��?k��,�/��۠X@ά�"a�/���� p;������������r����n������H�/c�i�*h�� -z��Pύ\�n0�6�^�ؘ�������ȏn�&��F7����2ɘ3��ad��2l"��ݒ,W����p�n�/cA�I�I��	�;�NջM�ؒ'��b�kO�n�fh��K�'�l���61�n3���v%k�@R%�(�X��OL����i"��s�� �i�Ѓ�'�[�B�n>�R�1�C�����o�tV��{$n��OpX4�w����}QG�'w8I�ke�f�|�RtI�4x`�T�T�h�.�	��z�Ƈ�A��bV�/Z��|���?<.�F�p�Y"���\v��Rj�:ܷ�_v	5V��W涷����vC�>�_���^Y�w�U �o��4� ��м�1xM�M[p�12�:��fQ�ҫ?!C0�$.�q��J,Q��D[4e��$��(&�.{�5x���&c��?:�K5�.�2y��������h>͛�yM�!�TMZ��~a����p���s���� \�4:�{��q,d�ft�k�T(99����LM�ߔ�w������M��col�S��g;{�Y�3��﹙�W��}�[�f�����n{����Q�M��=g��C�ȶ��v��	C�lՑ��PH1B���c��������i�δ #1�����i�� 3	!>ࢻ!ZrfA���?�$p�榨R�P����^�{�8j���6��#�����ޭ�={V��S�H�#u��g&���&��,�G����Y�$j�
����0rytPP<:]P���_6�{a��DD��T==l���^�)sS���d�f��o=���R`\��	�j�YK�
nZ�Ðr;���&��/}�L�8خ㯷���p}�5��v&�1k��>�W���Me��	.�q��Wfy?��m(�<��y��\��+�׽9g��HD.|��#K�v����Ӽ"�$��@�Zq��:FIP���gj������d���y�͠����l�$�����I�3z0H�C��pyl?a� ��7�Z�SH|�E����6>>��b�"�p�-�N���o���=�9�^Ŧ��͗񐝝}p3�� �� k�����C�tU	J9dr�	s6�_�� �2����!�QrX�`$��P�gGF�z}q�Y��	Gۅ0�EF������m����7J�"��1�g�J�-S6�Ǘ����/ҍB}z�~��%�����5aE�����Fc\�3"���r�?�Wc���i0s�;��G��Qg�8NI��="P&�
�K7�]���s�5c�=�+�������&��-�
��2��z�}�i��ג(�d�Z��e�u�d�;��L��H���%yn<�����������C����Sk�sw��K��=�G'�bĤ�ea��N�nY4�`2a��͏����ebJ;����Yѫ�+�z��_~y�OTm��h�w�jҴ\9� B�)P=C|�
T���o6`(\�!�+S�f���;AU��UgZl���&l0A�g�A&K���np}��V[@&�b�?�n��� � ���*�
�}��7��	3�V���^��=#��
[�"c�./��[�\"8�1U=c�I�4a�.�"��Z�uGPr��0�ʤQ�b~�;@�������2x�;�ɖ����������eeȭ]R�?�
:>Ӗw�.K��s��Fד��4���vl_;���%U}��m?J)Έ�S}�jU�"�R��$���uyl��g��27����'
G��e��/��ێ��$��ȱ��������"{^l`�m�ίuWz`��d-[-��3����b� K���<^J�jy�6�
��w���N@�����v�x�/u����#yٌEV�}7�FV�9��&�f���p����/�R*��٪1i-�;�P����4�}3h��KA�e�)�!���N��g�����'���e�;"RZ���s2�lJ�΋�3�.�
1�y��[�)F��fH�Daf2�1Ѧ��?"��Z���_����9�&�Z�:�Q����l��~�r���y��V�v�������m�T9�w�d8���ƽ��P剾���;������bp�������l����Q}��qp��>��c���j�����\�����u���2X�΃��,�Br�1uBY�0F(��< ��E�����o��LAq���{\+8F�5���GeЅ�X0Eww�TG�g�Ԝ�O�(��J���xY��D�wc!��H=�y���ڡīT2���t�+����>`�,I��D{�6$M���nN�/�Y��|��>!��"�4!ed��9u�B$ޤ�i]��]�A�x���u�=�1��Öǹ�c��Q�5pi4N=�X�=��b�8??v��w���$~��T��f~'�����������ֹVW�`�U�n���ȿG�^MA?m'�'��Iep��/u�X�6�!���gϋ8�*[�����|�OfeE��)7���?�2��F0N{����Mt{�_����܀h����'���_�f��yv�}Γ�<�M�N2A�(��w}HgJ��l	��C� �VZ.��}yS���Y�
%}r#|!�_�^�����i]�b��<�RL�UZ`���U��<�8͍�;nJgg��ʓhݢNX[j!Fџ:R3º^�L�CI�/���0GLf#N���������c���,�/��	����ck�췞+�a���_��Y6�]`^�����Zz�QHǰ��+�/�x[x^�`�b@Z�)�??u:��(�����)�[�
#����T�*��&��b�J�8T����`�{��E}w���q3,p3����Qͪbt�a�����f7�*̱��RW9���:�i�H{���+�X82^6P&/��^ �.p��;1��y�:��'��8��PvK��T�gT0񏴾SZ^r�b��W��ß�+&���Wd~L�?#�m�A?Ѫ������OOO[�Pb"syic�O�卲2z��կ�����m���b��̊�%���e�"�C���/�����L\���,���ަkg�rǓ�j�f�sI���޼�i.۔��g>�����>��`b78v;grl���Z;@����7kc���7��):��V���b^�U�h�JY�������k�o9���t"��]�=���/��<�:���4�睯�/[�j�k3�1�L���)zzN�=>)N)Vy��$��9]�8�P���ĤÔ�8(���m���d1on� m� E�8��
_��������@V��3e¢�[����0?�N�:�ݔB�4[F�0�]���"�"8w/�Qy"�}
0���q����bt�xR0i�`��S�4��Z�}0a������cK �L) Q�X�dq����� !���b6��l�z�f��v�3��B�6��l�#�~�s���g���w3v����5�x���)�O5WY��Ї�?��j1�Ȁ.��E`־j���V�[��x��h�`{���2��~<�12�$�U�=8Hsc�6H��W8e.��~����}*K]*S2�rcl�Z�Z�P���r�c���.�gV���d�V�p��a��	��.sn�q��0� 2݌:Vv����|�дv���C:�$jW��gX\K�Ij1(���%���CXU���H-�(<�ń>2rO��֥\�D߀�Z����w�v�ؒy�o��ZD�q����ʔwy=����X�r�<|�� Yzl5Q�T�){�Z�.�@ťc�Oxڤ�f'�x�f��^D���y��	Qx�Zm\��⬽��Z�A��+��xK�@	~XY�l0��CfX� �����o�����0�]<Ɂ��MT�D]������F�<>!��cH��_��1���Y����:�sA���虜x,�
a.�nb��6��fϽ�/IM����0��p%�&��d�d����1�giU���<N��L7��KdT�s/���d�Ǎ�_���bjY��8F�،���o�ɼ`�Bi`��~hly*�EF�dJ52__������^p8���X�>OZ�pZM|��DX�9��d���n9�j���d8���ώ{S8k�o��'��
e����4�,�ϾQ,���Ws�	��Q������]�O-���W���/��D���c�Wn.�E���b/zb/�ӡ�<�O�(�V����A3J���ဂ�nҐ|Gk�o�ˋD�]s&�|g�n�.�7�Ր/C|��,!ɀ��Hi���Հ�]SF�U0Ȟ�߮���`�d~!j���k��%VR9��j`��W��'T_��X8��>��'�
���w۵k�ym�Њ��Z^Yk�ٶC1c Ñ��r[�ʲt]+W�IīI�v���cZ�<K���w�}����a&^�:�|.�y�|���B5K��E���/l5i�k��m�=56�[�4�/�1$�a`A�Ef�6�x��Q���3qޞ։R0����'+D�O�L�6Fq2|�;��[�[��A�������o8Vŧ[�n@������`^��>����z�ʎ���{���e�C6A�"���$�)*~ְJ�q����(eRƟj�R�S98��dV!Yj����?
Es�����ȭ��NJ :��?�(��.`�O��X��?�����yم�c����o���]!����D'Y=Y,o{a��K0����4%&bbDy�������J6��$Gh����b!I�2���탰`֦~R6�҆��5��r�(��E����Z��xb���z�+�}��a�����}U���r-�#o>�פ7��Sy�s`�6ꔨ�^GA�v^��V�vBِ@���d��o����V��=/X�	`)��{���� j�> h�;\�6�XE�?��Ǒ�ɠ�I��ՙ�Yu�Z[M��ηes#�/�:����ҕ��F;�o�S^k���~\�s|�_���E�w-��Q�*��Q/����I����?��|G+��
�&ރ����d�(?�2�I*��J�<9��nJ9����<�����DtG�7�~�|c(�I.�N�ve��́W!��n}��ll���ܑ�$����"��������tM�e) C@ �@ր�Z:��Ӎ��,<G
�}P�$�MT]�6؄A3�������`������M.�8����L�z����i��&�I��ESn
U�a���gO��?�8ޑ+5��	nG�����k�+�C��#�,��Z6�Yk��5����!��[�Ϭu��Xlv�|K'5����a�+������D)�eG���[bߪ2v���R�K��̺B4�\0���E\�n�S�(r��kp����!���#���O�?r�_/"GH�k�LH,@�[��6���@Gz ��m�$FH�sf�w�����p�n�ۅ��Y��;�{,�׀����uȟ��;_8is�����!�e��U�p@�WM�>����ѿ��ܯS�I9����`oH � Nu�&��K}��))�Wr��~wE@GM��`m�1� �7L�k�F��+ԕ3����iF��K�=Z�������QV�5Q�G��;fR.`��0G<�-c��
�0;�?;��x��<�R���k��c���\�)�<Ղ*����K,���{�{� ��a3�!J��؇#����ݚ���Ex����$�.�����GI�Rf�F6P��bW���a�|�k��4�Wj@5ۿQ܀�����O�`��ԅ?��7l��Ь�9�u��썃4rơ��G1D���B`\>����[0Fɰ��.�:��
�=N�_l�	с�3^�6����|�Ĉxm0�x7-%P��Xϳ`�fʺ�S�˧���c�^3�MT�W�H�U��;�nׄ����1z���Io��l?��y)Y��8s���٪�݂�����=g�Gq=R����t��� �:,�O(Wf�q��W���S+\/�`�`�yF(�XW$cg �T��������YM�n����fAM��P�W����<|����
��v,l��6g"ᨅ�wt}���4H���Ϫ��Ȯ-$�����i��`Z��;X-�&CF�|�.]�X��cF�EU�gز�O�^ʹ���F����F �(r5�8$z��w��By�Ƕ:Ln�����_(��v��~z����/`�Q�����A��,�+�z`��ޣ�,,\�b�f(VN���A@�X�q�H��fo�{I�|jUW�h��ˠ�u.��OOP��?h�����DRF��hR�t\��r��4J�y+%q� S�yf��2h��7W߉�=�
�:s�n-o�cb��T�u��:�_}b�+��l�(�wcբ��ku��l�Π�?�k]'�|���%�F�����OcJc$#9~�PtK�L�a6�I�	G�N��"&�wh����\��&%�W(��cQΪ��R�_!���a�r�4ģ���Fec�^w����#����wl�W�Ze���U�(=���������/}����7�~��&��*,�&��n�W�D�U� 6����w(�Rd(�9���4����q�'�G�5ʐk�7��?��B��%}M$gͦ�n�׋mϨU���NI����&�Gz6�5��"|���i��Z�I�y��)�ʪ�Jᅲ�A�y�㴬d����!	�WK�~���<)�zt��o	r����G�]k�`Q>�|.�wJh2N@zM��41�o�_���w2֢L�zbV[\8�i���o-���|���#S-QE҃��{O���je�2Y[��ܶ.JR�U-�Ѯ�v�ϭm�cv��F�x޽�m)B��o _�����,�%5�;�oWi�[$���ۆ�"&��9m�E]d�������iG���NP}�0�
| &�4�U@�M��[�-n��k���\�S�����^ܡ�ww���)����{��\$�f��}f��4���{E!�+�QxM�q�-����n���;u@H=�=O��-�5�Jbbe}����[]��k-���U^w���f��Y�"䇆�8�~��~���Mƀ^��;��[��++�e&L����l�u�~+�����.�5P�����Ź�<��6:Hǃ
����v�*�G�z����f,R�|�ť��?_o�a�p��=Zc��t�Y�����K9��r�T��q�qƤ��]��D�c����$cDӒұ��E�H"v��X�ma��[��Q�ü��Xo�2��b@�>�s�͇�N��j4*S�YG�T�u��\�]!��%�ik���ꘙ����v&�k��J���ĎY�s�v��y���[ 4�#��.e�yM�k2F:��mS����@�"��4�n����i�υ�!|���Btp�ʂ8��8#� � ���*H�slA�Y�h$T������98���F�5�?��h�y�71���xNR�Т�����.P��>�v!�Md�Ż�ς�x�am����f��2����}�cU���|�^X��>k������CS�hlr(�"|�ߺ��$�IH�w?��v��(3&�d��H�����_���@��P�h�YO?[���UO��0k<c�)�*7�����и�bVJB���ͱe�tXry�ݷ�vuH�0h;S�lw�<�ҢC\�HXV����ى�����E�Z���	�P����ƞ�526q�K@a8��o�݋K���̌��E�y�!�ۗH_�T���E��'�yu�(-��a���Ri�p"��(�j����}2L���V�1/(of�fo9/�{�X4�SVB9��9Jf�Qv��W=��:se#.^>'[e��K��,����F��Vc�gea�ۘD�)�>F���5A����Q)��_%��Y� ���o���L�@+�m�
�Pr�ǚ�8z�jk+���5w�9���e�:Γ@dd-��o����Z����ާAcC�b'���CŶ��þ&�6�D_ĩ[�g�}���i��#ޱ92!.5Uk���Ʊ���;�����
|Y���H$GDaB�m|P��
D	��*�L.���N����S���%Z�t���$'�|�Xߤ�k�0����wPD?�p�Zՠ�8.1cQ�����>kk�!�����~��u�vl��$�z
(�,����w(�y������	j�
��~R�`p^�~�5�+p�����9bV�,�S]U�{ΒU�/`)砡�v�y�{V��F�<rE�gz�B7�V^��%� 1y�L��Ӵ�S�rf�_�� H��T���M�ǳ:�wpd7���\,W_;�*������!}X��J���Xk��*�~g�I�}Yߣ�|I�c�g�����{���LvL�t{���CE h.��k���G�4�Bb��R����G\��kX�f�z���n��gX���ɺt<�X�%ސ�es%������E��d�B��;Kh;�I�2Xn����.S��)e��W�?�c�|gPSٸ����؂�E�0�|Mz�?0�𷭯B8���R��F#�h'�*K�)� �~�j8�d;d���l�j1𧊜����}�~�7�k&�qe���zj��Ґ����Z#6!� [�HS��f�1Y}��e1�L2�>��pmeA�c���#cb�=H0#sƎ*;'�f�W�'�|}}�U^��֟a�> �Y�*���`���˝0�a"[htg�I�]����.!�z�;8���_@s��>Z]��7���onn�3��&�܂W���g`�����\��}]τ3��'¶5�(�$�,<��7����+w1$0���8U~� Ջ�����ek��Y��Ox�uC�{�` Q��%��ŷ�G��}M��{�jrLHM��A�*Fd��R'�Z�G��{Y��^�1hK�?OLn-1�� l�﨩�'��d"@=�F���_%�F��P��V�X<X��ͣ�LHk�,��)1Jq2<�G5��CHc��{��"?珏Y�-�^R�����Ez)*��>"���?��15��FH������1.l���zw��g�����׽i@}{J�fO�|ꩁ,�J�K��a|��Ƃ�"Y�
3�vx��������e�K��_��6o�^�7_S�fr!^�'<�~k�Ծ[�_���߄���'����IS���:,Nl���f��mw�� s�2Ѻ0��� ��k��,��˄[JfG0�; �c����u �Qy�WYJR7/�bہ�~W�
�3h�59{oV���m��O���Ơ��?�M�@?k�L7+;,����~���Z�����ߩ�m��Y��IEd�i�z�d���FYZ�`k�b����ɒX����a7�8�!��,"?��/r�,8�'t�O4:��*�H�Fi�M��I��v��{��dRn,��*"��gDG]W�al��Y�E�#\�P�06��1D��Z��*�J4��Z��դ��֋2�L��4��\�5��&ː�L%nc���d��Y�ڽV|l
n�A��]ϋ�E�e{��|�|����{/�O���#�?�����{�,f{�W��I�3����:�=|[�;��<�r\1\1�����d6��W�!�S�\��j5>��k�/���_�(�����-��UG���d���c�^c�i���.���ͦ��l�HǤ@�N�����+��6�l7ʧb���:oL���6�};.+Yؓa7v����I=���b�dJ��;_*��*ۻ��}��j�����YF{oI��*~%�.����V"1�Es:lWE��J.��%]�|FU�9�)�=�-ь 2��ڭ��l1��JbIf�"�  �u����]Ҩ��BC~�b���nzV���:s	��* ���h<J3������^)��F�9���bK�����R��e�PW	�@��:ZC2��ê�J���R�~ᓝ�-"������-�>���P�?=�;��8zk���V�����,JLĴzj���Ỏ+�DP��A!�W�+�W`��1y���˪�Nà-0�X~�Fn�l�_���=G�����G�E��x����ԷטW��킒����v�'^{�3f��ă�G�cA�j:$��sbQP�f����˧���}k�@��Q�pWN���w�a.��eu�;�g����X����5u7$)"M�CK��gKo\������uͭCYh��˘�$�\�3i6�C���~�BH<CͲ<���EJ�������w���������q��Ig'd2Z&����_�)G�&���5�mm��|_���w������|ta�6����t-޶�S��g��g����9��YB�-\�q9�s��z�9l���ِ�2r�CS)�~�v���吐������G����l#�7��}�0����(cZ���;<\���X'"��G�z]��f�|���2K�i�^b�~\�0r(U4��_��x�Z�n�Ʋ-��o������Q�]���f���ȍߤ��6{��b��k0�[�8
��2��ʨ
{l��QGk����NW��{d��
��u��y��&1p޷s���77O�ӻ�~�����)����D��L��.ೞҋ���U�
�NDxվ�C���f�fW�5W�ӛ����Y�qp�w	`ǎ�� ��(L�L=vr�<�ii����|�<v��&�}0�l�a��q"HK���T�����.F����c�l`~+[/��3������<�>Ffn�g-�z6�8%�m�=
=U��~n�З,��7]���@�`�_1P�B�d���R)	����|}$Ն��(VC2�^s��J>�5��}o�Ȟ�c���KS�l�f��#����#m�#�����	)���Ǯm؏duBJ�p	��^�F��̷��q�4�2�2=>�g=�E�>N�vTƿ���9�>{x��w�I=H	�<{�7ʟ�m1�Y-�ܡ�ҭp�k��*_(�ɫ��g�J���#�r��қ�}[�?�9��	H��Σ�=t��0J`T�܉~"�����8��HI��ޓ����1�W��?����z�}P�-�W�=d}�"��5ynNr�Ul��׎0�]�{�����Ph���bw�1i�n���U�޸*^qe(��5_����׫�Qf����T_�oC�E`CL��xcw����x�����\,¥̽c��*#�L�ĸM�iNY�4z_���	#�hi�~`o�p;�[P��[��5�B5��/9jD�l�zI� T��[$+�;��n[�C73����$���t�0I���ޤx���]Sm�ּ +��l�'YD���3���'����8SH�:���:Қst���HA����vߵ�����}[7�F���g4�͋��1� �������+#�-���>Wҷ֡�EF�l}i�X�Dv�њ���Ob�΄�&2��a}���߲ˇ6h�-���7��H�kL�R(��C�T�b6�
]/����!�I�,�^�fVe�K�����E�۫sze>Da��o̿Zʧ����/P^����1g;]�/��t�s�>�/�������Lg�[�I�^�po����?�;�¨P��1�����ХbHL���]���Ạ͒w�k򅨟MW�h�ā�d�ؐ{ִ���Y�o�CH��I�*+c��Wqzr$i�}3l_���wrv��X��>x�3�6-��2.�%I�d�i������������[;���R��;�/������2�����>\_�W�[*���S�?� OH�%��w�g��>˘S�<}�+v�y�9��J@�ڿĞ�s{�u�V�ׯ�0��<���ڂ�E�bl�ao��QJ�u�5�,��$���$�,�O����&Λ���;��'�i�l�&���`�J$*�d��RJj���A,�k,\=`�����yf�2~EzF���-rE�{ɪӨ`����h�7R��Ib��ag� �a�0����%�3�њ��+'[O�	�L��T[�����뙪c�M=ا}���O�^i Id����6�Vg�_�l�1����bsM�=�r��OG�F/
�5-�����UcAm�c}��H�l�kB`߭��T��|���!�sxM��7b��%��_�)o_s�4[�n#�И[��5��*�g��b�tg�G���Fs��?�U��S���/�j�eq��(sz���0�\�>S;���D�,>�B�� ��>�D)��N�W�2W_�C�c�Rx��驞��(�)�Y�w+��Z�_e\Ѧ9�Bt�e#���/�0e���|^M��w���n���Lz-����X`�4�X*;���ehl���?� 2� sn�0��}᯵CÂ������j�Ȏ��B�!vA��$���?�F5ij� 
'V8l^jC��x@�!�Q�Z��Ĭ5I\���8�0k5@�閳��f55�\^{q�G��֢�"��}}�I=��]&K�i��������/fl�3R�Flz��اXs�r�YUv�l��4�� �:�H��.>TkF�������䤡=Ǧ��£���?�!���q�k�"����	�aՂU��4�m|W3S62'���k�[���-�+{�����7�([���V�8��������媮�T��#�����.��Ύ]H�)�ۮ��m��\�I�O�ѕ@��J����<u��Sd~^^@�	��X�<c�#�HjM�+�D!�$~�� 3������y�)E?v�`��>������+�r%���f�ϵM?� �R����v����xM.WԮy�bRB�Bk�0��-#,տ�hB䘊y�q	��eX������R����E��e�H�m.�ŋo!���3�(���*���yc�B���\s���h�'�p���2b+����mo���U[�gIQQ�0�BJ�����a��Ns�8�{�i/�.�;��^)-��(|Q�q�&وG[?1x�o�{��w�V�9��7�1s�k��,���V/K��(�n�� M��,V���7� Ǒ�M��(b���>i�!h�\|�};���܋� {{���~4HC��Q �?;&hD�o��dP�&�-�2�,}*��@�K8_�7k���{Mv�]f������i]@C�ay����Z���zw�i+Z����� �\3I�1I�x�
��� L����I�a��b�$���+Z��"�E��ER�;�寶�b()!x{��S:�K�H�l@H4*��]�G)�����'���}���^�֟D���GnQDU��ԯ?�\]�y���6st��W0(����Sz?��7�d������uS�}ar���똤�(��a�A�^�Wp�L�\��n��Og���,=J`�.n���Q�����s�c��! 
�URr��M���&yt��#V�N6RMge�A���IC���5�0݂;(�T�U[s����^cb��c�W�f���d��QKJ�pŔ���#-.RB�D����aA�b��uR����U�,[��_�s�h!����7�(�$a���<xv
/�Z{�����r��r�I��*��b��0e���C����q^��?j�Z���[�~d�kV�7y����9�ӏy�u��e(3}.z@�IȂl�n�vE���& �3$����(y�IF�M�6�j��(�9N�/w�	a�o!MY1=ҰVA�Hٱ��?�t�6.��^%ћstZ%ibBao�TKWs�a_?��F����m��M�V�"v l?�X���B���p�����"�b�������- -t��/���9c�ƈ�NI�Ah^������F���PV��ЎM�d�����è�7Y���Wg$:4su�T����F���x 7��؄�n�5Z�zi}-f�Ĥ��LyM__�ҕuW����v)�?Mġ�(�5D%�OD��w1m�8��͍A*u�{��׭����]�gj�� �]�t�n����
=���A,���<�v����Ni�_mP��#�^L�9Gc��*l�]5>��4z["G�8q���`-��֟pm��"sՐfj�����$��ܞ�F��&�'X?����CC�ye��In��o?��盧U-w���<�ԣ%([T~�L��USf�aw,�їΕ&�ňp��e{��?o�����{��S���5Y�~�a�Z�P�&��� ��t	��Y������b�n���у`�����SS�;��&��hеD�����T����
̏��"��N�#T���D3�O\>�nq�&D�(�M��&�h��
���ҳD��kWZ8�P�|F��q�����pE���f�_�C]�)lpf�#����\�
����z�˿�-��2k����)�*�Vo� ��5�ps P�����A-Z�~�5��R�z��uZ�EOs�e�d޿����lh��O�QI2ɱTk�@�M�Ã��?V|<�	wt�d]�6u��`2���u�4g�Fy&!!N7�ig��^�� Ϫ��t��NAb���Һ� ��WZ� bﱇw.�K����Þo���Y@���_�}ćy��Լ���%�]��
	�;b���G_�?/X&�SeG�8�:W�9'�s�[H,�M��N?������P�k�F��|�P>���h�;��C$����ɓ>crڽ4	,�v+��z.j��!xݸ�{�yz�&��-���x��VRB�y��#֋M��(�P���Ske�b��ݘ��x�׏.hik�RdV��h��T�������Dݣ�i>d�[�\Jd8M�H$ړ�6���9a-6D\v��VKj�,.�7{G�ѻ�}
�A�;��ݢU'��4)��OX�KeK6��@��oQ�q.�ޮI��~����l���l_��T�-�O*z�I���߭�#���A@=���2xe'X8����#��k�E(Y�iL�SY��Ψ��9��"�x@���&`h ��8�B�Yu�W���L���9�߫a.b�Y�c�B.hYX0i4�d�X�Kz�s����;7=����iH<���=x�/�	�q�r�����D#7l_>���/���v�)�=�;;�������2ஶ�P��a���X�.آ����i�6��ǳfSV0�)�)�)m2H�u���NT���� �XqG�h�,�0���	s�Y~��7�Z�%6�h���X=����μo�����SuL�,�:b	NWm�����i휫���N�u�;+,��;�W\���'�n���������HM%PBZpH[��s 
	
�@��R� _sf-9�u#og:��5؜��f�[y!^�;�<��y.H�uKK,��6��j�L��v���0�&@����&k��g�gf�H*��A/�^�w��~�s�J�g{�Z\AJ־�Ɔ��[�ob�?���\4)iZ䉧b%��%�Q���A��Ņ��N�YG�4�Gg�#7:�
��N�j�M�Q���f���o�n�?�)��XD
j�nӘ��}��/Y�l��Vt��%@����o��0^|P� 9yy�k��D����Q���ӌ=-"+(�)������z_"Qn��''�	�a$�Ю���w���b!���K���k�s���$�V�J��5��<6>14�D�Ρ�~/GD<��!h\���..S�@%RPq�9e��5��f/}ǉ'8$��a. V��$����7�l�s�w�M��1"`���0�{���wdpi�P��^[��!�憗
���>?G���~����nafȪ؞������?d�
�q���%/�;��`�Y.�B��g��M`���,�Ih������%�|�7�֑��rB9; ���9���w�7q�inp�o!���u@�b-#_�d�%\C�'��P{��m���=��s���}h��DUӌ��&Wѵ���_�Ż���np8�J.���3��.�٧{��8Ӣ���<���2�9�CnQeشاdR{�-Q���P)�Ή�*aJ�h!�0����S
�lM�l�WA��6���}�|xՅ� �"n���'/�s��x�+��e)vIO6���M�v���� �.�,����=��M�j���
���]N^��E�/�\<w�Yv���t�R~� s ��OH`u;B"����0V���1���.6�����F�<�d� Z�|�9I���j���G= �(��Q������0t��[�����42/s�]�l�5����<�]~��zMv%���b#-�%u�:���s�fgUj#�u)�w;9�#ܭ^��J#c&�dٮ�#Q�m�f�~�}�G���J4C��ouԮu/e��E�Ŭ"�Os}��c��_�KR;�<�+�)U�A>H�,_..����ihB���XQ�Y���+"h% :Zp��ʇm	�8Sl�HpS��t�ܧ��U��$�ȈT@�Zp@z\TY�,F[�K�/�	���4��|n|[8�>|����8��l�YJ�*�����rsk ��©y O2�u+���t^��O���w;q�H�f�.E[���3����etGI��o�!0��M����L>jrPC��-su����5V����"b�[�,���L��9�('L_6��:پ���N�/2'P�Q�Pus�Q�$O�s<��|:f�3ۯ����[�����"���ץ�*�,  ��o���S�����w�
DB
�؆��iм��=cW�ؒ��V�hc����6�{��DmP�z$��=ӻac"��C�"-m�+SSS�~�[��511qV`KH����C|��p�/
cW����X���KBZ��e	�>o2���cE<�[�+p�&��"W��qI�v/�����8��7}U��aE�r����c/)k�ٻM�4Y.;6A1�Xc_�X���/W��vj���WBoȟH���U�U	����M����>�h�����b�&�*���E�{�fbJW�Zr�(�An,@�O��G���6=���_g�ٞ�1�]�ĊobEvp�e�P�YZ�zNbo�1w�U���2�����V�Z��m�6Q�G���,G�K��ݳ�C�I�)]P�^�s�1����ȝ�+PR!��ߕ|-�-���,;=f�I�>ѥ�@�A��t�1��
���1�&t��t\��Loc��.3���8���=�H�*����dIu�^���~<�\toz�콵ۭm�#��z�(#�)�x�w]�2fVg����pY�Q�nՄ.�=���^�i���A�V����S��@�� ]�������o *#l�
U&h:]��w����8����!Q�6P����F������}��������@���Ҕ����ԏ��pڍ��xp@�
w��D�nP!�>#;���J�|�ݖ��4��!vrҁl�!���C��"���q�ĳgjhI�(#F���^�hr�L�9P��,UN�IC�b��eI.�R���m2e�P����a5�Y���B�����ٺ���S.���CC�zz�7�q
E�����b��O/_�Z�n�k��L321m�0�(!4����{��ѷUet`���*}3�P����;�@������'Q�0����w-��۳mU�� ���{�Ѝ�2g����}]؞�S���������C��m�O0�і������� �`���N/C�hl��K��\ tp&��S����:۝��B$��N�~�{�8�����{b�����F��h�-'?�s ����EP�/����Ӡ"���z�wj�+G�po@ˑ�� �~�7>1`�ۇ�k�]]�����5��9�Y�G���<��2�f�����8��2��M�-rp�:f�W���f�S5ꧫ��ul���ռ[W�2���h��'Fe= f��'nqZlGǸ�Do}����	�hR�	B����I� ��ᮮw^w'F��Y������ɚ)s�5a:��ή]cE�U���=s�ҟ�)HhV���Y��fg��S�*(��r%Ȥ�1��$�/y6�����'ⰵ@�a�?2���3����}�]'q6�)�i����g_iE�_3�i�Ś�}�G�%Ô���Y����_�`��[��X�����?M��ZxL�=�Q˳�V�/�&���?�]��@��5a�o*�C�L�,��cD��c��Y̫����t���$���M����@�:
�U�����wAb���=�n�["b=�|^^�1����M���[��e�K�=�@�^+��%�]�+�"t�y��_7��lxL#F+��!ÛS�-5��O~&%+����_�S�QK���9ӂ����d��)bCk���IF��&�����b+���\�o%Z���/{�f�{��77�G��-Vxѐk� Q2{���j�.�U�?_?��w����SI��I�C��b� ������d`O2����3Wq(��Gz�Q�櫤�w�ǍK�x��+��[6����s3z��8J���iij�cp�4��o�GZ�R�3_%�;i����}.��u�\��;���wm��\�\@��R:�&�z���;vխ^��������^�^��٩�p�3�a��jn��� ����Q�����dB\" �v�x}�_kk���q���[��W&]z6Y@t�R�53�c�.��Q�Ynv`�f���V�}ϔ��YY�ǧ��n�n����;%�]l4;ތ����U��ge�ą�y��w��)*R$�c"��5k���Q�.�~�r�u�ҶH��(�B��Ʉe�"?7^���I2kxKjx�E�~R!�[��T���z�>+C��e�v�)�*g^�g���?-��,�W�u��øn#����I�^�w�/B�{��a�>$T��li�Ti�R?&1Ds'��"癿:�k6����]2KIo;C^�Xs�)�����hv׸�L�9I���0�h�Kƥ�n�4%���hp��(���~�C�� ;c�r�j��
��S����W�<�s����ī��{=�"93)�F�1���i��#��!�Q��Q't]i�G��k�7-�+5���S��F����v�/P㣽˜J������龣���*-�����ӳ�Y~�E.^�	�8��bk�Jx�x[kv��<A�Ro��l$x�[XT�.�������:)6���Ӟج�mօ�>)�a��k8�69BS���Cf��*��ʩ�֘� �z${(���k���SA��6��v��k,�Œ����~�F�qΙ�:q�-��ͺ�����v�'%���]ur��d����k��y�[ި�<���8˛_E0����q
�L�ۃaqrc��)���
�.G��n��ظZ��^_�ϣ:%���^���U2F�H�..a�p}�FJv�0� �(1B��S�r_m��%>�����:;Z��J%פ3��B,��ӭ!�ȦM�2��{iIugZ\�3�B ЄJ�^�:�d�D��gl���P9��]k�n-D����I���\��N����g�n���(��tD���WX��%J#Vk�ԝ��������.����c�\�A<x���Ӯ�);�)A���$u�9��%�q!Ef�D��;ձ@�-1W�l�k�䚡��I�7���G��e,i*���0G�L��x9p-���m5�s����r%��,a5
S��a��a�#+��4��8�d���l�y��/3�J��X9��@(I�^�����V�BN<�M�9�X����e���E9�n=;(cA�;C�'���5)�y1��ˬrtd�9t��V�������I�����钜��YYfcT�*&�S��.��R�Z����?��	=�vi\ R�xz�<���`Wk&�T�������W�cj����ӓ�^�Eo�+R�"A�	�� ��d���=�~�ǔ_D�)H�[��)N<P�q���%��+wȰy��ygs���DG��O���.��R�DgG�W�ci�`��=r$?���"7e�B�|EF���� ^y&�BF^l�b�C:h�&*�.�:&tQ%�D��vB���Օ{�"#���$�����#�"h�QGUd�6��)��9�%M)J����7�4�z���w��X�GZ�����p9^�1T)�:�<���GAn�_�Lֿ�sr^6r;��Tu����EO�7��-W�~�5�8J��kvM���7�	8����X�}�~�
�v;;�a��f	\�d��hDvn�XN@]r�����!;
J� ���1Q�����S�c9�DŖ�Y8�U����L���Htឰ+���tU� �h�E af$�l��#KM���&qǓ�T�!�qt����0m/i���3bP�@%_��Ҫ�4>ν],����JU�g��-��hŁ �����������z��ʌ���l��P��8B�ס;1Z�=�W�H�}�ّ��9G�=t}-NC
���Wc_�w�7�������>"�ow����_l��l&���h����r��4P��p��X���,��\q,��-�x-�q�b��B˯R���H�M	P�B�<)f���2��KA��I�{��j�8�� #y��t%�b���W�S����%kt}H��'������lu;+Ԥu<�+�)�'�#�� �(�䌂��-f�췘O���--���N�yU��b6�l�FC�n�����.a�j]Hq
�ǷoG_e�5��\_�ؙ���|�܆�b��,Ý��:ѧx9j(�C'�Sb�漭P]i��qT$S��SB���5w�A�M���[��+ ����9�@�$2����x���&������L�O�=��5 '�pÛV�t��300pp �T���BX��|f�	"��v���8i�6�ܯ�b����Ey�F7�a��c:��ޑ
�y����<~`X���D�0�l����Z����p{��k�oD��j|EI41���S��M�Y�Opw�����.J���"{��ִIE��gl$�����l��hze�w�`x����1�*���40���敏ф��HF�u�g#�S�����
���.����<�䮱�1����B@ڶ+�\ Ʀbj5����j��}�٫d��\�\�&6T�I������bj�B�D���Wo�G ��7�]ܽ��-��ܟD��x[B�B>����M�$Y3�J�oRH1}qx��`�����**عżt
ۺ�f~{|���=�d�C{��b4�J4�YsA�_N"k݅��п��	";6`�ֿ��D8��s���S�F��0eI�z�v+���w��i��� ;3�{���u��*ۡ�|�<���7'V_����9]�!�WA�Z��� ֱah-��ǫ�-�`w?xb��&��Qh����{.r����YH3<�:���hZ� ��	-��؛ur�T�����X�8ю.h�aI��~
6ٔ�I���4�����H�I�.i���E�J��F�3�c �����_Q�~�_�qDċ�vvN�A�t��B�S���� �is�i,�#/��#����Y�����n�gO�yʼ||�Yi���������Є�����	�; >��Rf���<�L��۷=nn�zw��B����>3���p�P��@N�+U�!(-ͅVO�M ��&C�.�9�6y4P����/555��2��_Bn���5	�Vvv̠��y��s��QŦ�q#򋄀���_�g|�	�`��
�����[�,�s���?�@c����݄�^r,K�^�����y�k��5⒵?���x�p�sO���%�N/M������H�X:PÉ	ź?s��4.����Gv1��e�.�'���e�kL�g��ZfTL �=�m�>��$��t�f,j�L�Z��(���$q�ibN³[�1@r���uG���帹%a9GOAA��8�������Ļ������Q����˔�L�L��# T�V�`~u(�b�ܴ%:�ؠ�W~�V\xOu�	e~����ͫӛW�5Zzgg�饹~��_���&�+-�和$7��~���1~�F�{f�vQ`l�߇�I P^J�ׁ߹@�~d���	����*>D����}��7��H�m�����dy���|q��+�a��.܃a*�|b�;;�.%��G\A?��˰����*A��|:O��n�5����g��E�Ee�a���T�E�ۤ�����)���h�)��zq�@��<�5��9x���k�:N���(<˺�珩�7�����h�R ,�K��^K^���Y�h��5ӷ6iF3�@JR�6�}GL�QJ�}"964)�����=A������锯�j�U��3ѳ�Sy��e��� >��:X�Ϊ��n���G�H8�*�����ck.����|��h��Y�1<����ųFJ:�X�LOc^]�q����G��������z��A���ց0�O�Iz͢�ɀ��1=Yʇ�]���o,_>�M�����5CQE��9j�AO�ƅBV��i�^��`������O���MJ��"��\dL�!`�"5+�x�[���P�~<�1�<̜+�����*�+?a�7*�(U����]�)d��Dh	��:�����*e�c��|�|K�ډɶZ��	��L
�ɜ6R#����6_�3;�.���T���s�oBs�^ygTN���L�U�o��&�3�l���x��MU�76�-�4�X��\%Ì6L#�Ң�E?��)�O{���`�3��3&1q����W�;Z��D������3�Dʓ�`�=4R�w�Jl�v:�ʀq'=1.��:�yf�	lf����<�����*½Kw�l�8���6;XP�����o�8��t�^_-u���N����U�<T.�v|	-�fe�-����Pr�
q^���z&��/83�W�W�)6�66&{��@�������Ϯt:ot2��P��"|�n/�^��w�_�ޢ6�auCsf�`��>�'��T������6�gMa0}k�&���_�q��k��U#��hY8]E1=3����x���~��e�O�2b�9�g��������sH����p����xY�<\��뽽��^�� �9��08��� ƨ��R*��P�1C�0��%��sHU���R*�>��}|<�t\�~M�\��Mo��xP%�~O����G����#q�<�@�Ž#�*G)����飹V���j�_����fR"��K�J��Ƈ��*V�΂��&�H[�=����܅v���>̝h���TX����wo5tp��	l�un�a�YE͢�'��v���S@�$����m��p'��T�^��	���%{=.�4���Ϊxd`P�$�$5�e�|�zީ/��F�ge�������M�7�L���T[��7�% ����1>�BTR�"C�՗�˂A��|�f�"���!��W�ON���'_-�c�P�5ݛ,��p�>\]��V;K�2Sز~x�潦jH�.��S�8����E�*�2�ԯ�%��:��N�w��k�x/���!�Yl�բ�'��$a��G���x��4�����L<S�oH�J׳�~�	�cu�R��?�R��+4���:��`��-��(ŝ��V�ݽ��{[�ݭ+��/�4���C�p�������s��ٙ߳3�,l5:w��u6���۪Dὃ�Z1X4�����n���5�-�m�	{���6	�,v�)ly��un��^ZyP�x
wE�|M��=�X��4��ض����_�.�)�*��� j\!{�^�e�v��+�Ze�i���'�6>����܉;sp]��ED�z|��{���t&a��z�y� N������5� OZSI㮳�g�)J6u7�t� z"�d�f�O,�	w=�����$.4fN�����F��-ח�e��l�A*���+�:��@� ��K�L��O�i��Λ*z���	'��Z�gd&�	��jR.
���F���0�'��h�;�Z�� �1�|�?U�fX9=~�չI@��a�����ww���K��|^G�a��#KKB�=���=�.Cx�>��{-�\��$*���%�%9�]Ay�&4*��[L[c�͊D˷!�������w�f�����3�Y(��+�exъSs��w���q�����	�_.b��W5�-{�댩Յ�o��a#2�Ͱ�pՉT&U����)�2�.�Z>A��t�l����Kt������r��'��еB[�h����k� 'HXf���rIUM`���b�'�N�b����B�8�����,�!��K�#"SM;�����V�H��:�whe�P���I�7=�N�b�t�|�$C���J���/���z��p�*y�?kF�R��˽����`~"��&/�Tþ��R����`��̘'�����������s~���@�t�ׯ_�
�WoٕܥR̲i���j%+�̓�0�t��G��(vhð�M�W���Ձ#�	lfj��?�d���_o<��n���)o���^:�|&�Z���<m��lXؗ��~��^�F���*m�^�v��jn۶s�u`�� �������\t?�{;�ʕ|���_����Z �X>Dg���?B7�����*�ɣ+�۟����뾤�>�*��ݷ���R,�\J+w�8���|ݍ���0�����P���BHI� ��ݧ=%���ͽo�������Ib�Ruf�6��4bS������,�3P�����o�Uj�������;i��Փ`޿c�
LV�cV�D�U/ƭ���k��c̖���:����a$0rͰMd~�P�ٵ��k��|76��|n� ��~��H>J�):�t�6���ӳ�m��F���Z�Ǌ1!�Qغ��3�y���޽ޑ�"r:��Z�%��d��_^N�6Ŕ��-�ݞ0ԭ���a�d�ZY `�� C���w�1�59&��[���w�li�O�c����(��V�E��,Eu&�aIʤ��9�#a v�8Io���I!m��m���ahӈ�!<U�*�av�Ω"�C?f0�IiMX�~k�1��<3z��|	��z�b���E����r�_b�~	A�ǚw�W�U(�,Զ���5�!�2��2 sRk�X��8-S�0L�p}@��
���r��s��z�˰������O�5��z+���Ã����Ġ}�{��~�ݺw���/�,�y���䱣$'�{?K'�gm�=�$������I���k�f���_�I�?�|��T�/F/�a<x�&1X7�͏C��i�ҦL_Z&�zן����-��-�;x��2Jԣi%���`Q��ٞ��Z���$Dr��(|6u��>�·}�x�o/����S������k���0���<�7TV��Z�}8}8��y����*�/�;��uU��|9�T �`�|�N�}�����1�aIBS�;]b~7���s9�oT�	��"���F9��(3iB�7���'F���4���cR0����{���ЬP���G)�"��ǣ>�V�Z}`��:�cB����`������\���N,-;w�ӂ�.�444`�ˣw&T�#n�ɸ��8p+L�Ζ]�#Ŏ�gȳX,fD����ǒ$�Q��+�yJ�'+ϰE2m��� �U�PQ15n���0�82�j������U=�yH5��Q��h�'+a%����,g(���hJ-�O��*��~:��*"��l))򌞅�01q=v�hkz��Lv�^��_v���/l����,Тϡ�&B�);�>�#x�Ek�k� �A�=$�SB��X����#Q3�s���,=�E
�h��}1Ja*%~|�7H"���K�UWQV�Y���σU^�!L(o����#U��.�c�;�^�g�-�l�4���g0��~&�żm{E�)�r���Bƭb
��"ə��i�< bC�L¬�v5����=U��������r�bW��&�J�U9$��d��Ȳrʗ�����wXcn6;��k����5uX4���c)T���Z�Y9��mt�7z�h�Ҹ\�/��~q��ǳE����B�~�J){�	a�%nK��P���>�$��)qӴs��/K=O���&��l�(��z9,Z��}��]_��i�ɤ�5����Yp.���W.��bq�)�q�՝��K�*��[���{~@���j��bqJ��{)g�(t[�BD6��x�ٔ�.��ԇ-���Q�s}�F��?�zڰ-(�^1]�o@�䙰\3�k7Ŋ�i�Y������s�aG��XkE��5��2�@�G9@���h�+!*�w��i;�4u��YA�@������չ�DP�趋f!���BG!19)�����
�(�����]R����W�����_��#,����2���!b��a�o�VC���*i��S_�>]�K�%�i�{���r+k%1 ������%G���mG_IT�������_����l�U�'���?!�G|^\�'=�9NTq���X���7(���d�r�O0#�
40��Ze�I;k�x[�-�4�[������ᣮ@*�ǪU�A|� lqN�T���p !I�Bo�+��8�Ck�^�Z��i�"�II[QHK����b�,�6��Vt�/�d5��X���V����-o�c��w�æf�C�|^[�ǛXu�4v���Bl�4i��޸��|?����x׵5S��Vz�_��)���tTK�Y��C��R��j�M��6]SY�wPeAR���B��OH$W_�I}��G�r�1��^��x��(� �q����_��+����B�����k�$Sj������={!�p�I���R��v�����Xҥ�M���.N�+�r��SF�V�b�S�N�4�s+�X�n�V��Q� �C�+*<�����p�=�3��B��U��I�T$�B*.��_[a@�2�F���wr"AwX�}���n~J�Z<Y�
'}^�r��n�ȃ�AJ�$��2mI�H᱑�W��r�Gq1O���������%B�,�r����F�Ph��t��p��{����m��%L
��� n-�,,����B��CB8�e�]�����M��@�<��?fT���qJ�+]6�E^�tn�_�Լؒ������O�	�Z� s�٬WTRR�Ԅ���/��
�W�N�~�j���|�|K*�0��%X7���R� ��Q�Z=+[�*N!�:�it�H���x��x�۪͚`h�R��C�)0l�o�S�d�3���q�ruj��!ˬz��H�ztR6G"��f�nfN�����m��&�uu� Q�`�瑠K��>��Ik�� [��9o�%�ߣ����i����S��a�D�st���ތGޯ�9�͇J��?�ss��vȚyF�Fcʱ�DF�6�!�?M!�B�G�q�7���ct�3KŴ9�$�Ł�%V�[/mD�e�9��'�*'r*o����Z�w���<*���*�q}�#[����|q\L���5�S�IIF�?y�i
3��v�Ђ^���!̫�1�����U��n<F1�Cm޶����>�7��L��!��E�D�u�9�G��󐌏
�39�I~�1���bX�� ���G���K��T�p���& ��q��?�0Y��^3�N�-۹ޝ!�vv8�T�������8L��~i�t�4D!���l��n����|�uE6E� -r�*+��}|�ht�Á9�!ԣ���1x�UB�v���n,�u��Oh�򥰐B�_�8E�l�ݗ3M��T����!��›���H�E\��jG�"p7a!K�^Z��pR�{qN�b�!�$�X�R0����9���p�J��71��s�q�תz���$]��A��s�u�8�����뺚��1�w��*�l�ܠ,�]Bb�h�*e�.�č�oHd��Ӏ��Q٧��������9�=ʸ�ĸ�<����)om��:�����c���{�}�q�#{�%��D
z]�N�9�(�`��2km�%�Ŧ���vv1������EҦC�-�ѿ����̢F�s�1��wg��wХ�E��Ka�wt�6�i����69�W���?��`����=uA;NkyR�jW*4%�vsxtQ�cߚsI�S�2���UX�i�ž��\vt�^����D���dR���|-H�7�Dy�ȄG��1K����3x>���ۜ�_��b��C��M\�􌅯�h�R("ʪ�G��R������"ْĈT�4�q�w�`���w�M>,�*i�2K/�ȸ:e��\�l�����B�1�
Ш�N�<���1�Հq����V���Kj-HZt��'[�O�Qj9ZjI��f@�D�q�NK���Ô"m�θ�ж�� ����ϭҁ�:i�mxs�k�DƱVE���!#���"�v�(����N᠍�eL�w��>	�<܄�b�	h���~ʄ�M�>�d��Z3��+.����<g|z���$c��PH��N�E����&@�������l�C�� �;��I$l�����>��M��h7�<^�le8|׉�6ob��RF�΁:��*���>��H��ѿ�փq�t%Ё��l��i�|�(�ܙ�*j�'M�	84�F��FL~�J��Y�q%67w��80F�.��@�)��hC�2��`l0pd=���=���lϦ$@�{��z���\mH"�`ץ��!s�e��\�%g�F�f�c�x�߱14��y�M�{��~Y��ɿ��냊��љ�C_B��;�!��{w"��4�Tp{��1�ŉ���Z��}���]���������s	�hh��%��Q=�"�ykwոp���t�D)��T%�n�+�&�l� �z2?����k�D��)��.��O�j���u��5�<�������P���|IT/�-����y,��x@f���������|NH��W���J��vy�[f�W�@�p��E�"G~�]�E�֌�����.�%)]��}#m�Ba"/�^�)�@�Oc��Ë�Y	G*ϡ��>�۩qȹ���H��b�hP���5�7��:��T�F�6�g,�wT�rn����Rpn?���|:m۔�����5I���Z�N�Dh賉(�?���J&�e�zo��bl��Ft������d?wD�?tG�qS2� ��v"��~F>m��k�=un!��[r����߾=�G���4C9]q8l��X�E�(}Rv���BL�~2���|هK��!�8?��_g��=bi}����ԃ�`�X��ĭ>��||D�x�>���ztZqZ�h)�}�Ź��2�\���Q��-�iZ��i��t�s����i�2�J�8®h"�DІ''U>�0/�S�������9[�#?m�w4�6�W,#���c�k#��V�����R[��/���x�h�>�Sg7K����P#~L0j�z�Tx,DE|���u�"M!�W"�1��+$"ڿ=L�0��jA$[R�����c|��?�5cn%�d6�eV�aJ��Tx_c�]TH؈���w�Q���5n� �)���\(��'ز�� ���	�I"�>�!��Q��V<�Hu�=tX�y��~G��u��^_���:���j�!Q�9��8_(���D�u�!-Z�S��׵_,�:RD��KZ�S\q��t$&&��S�?1��PG�[TO�cሢPfQJ̒�G�^ϜJ F>��V(�D6��%�Y��=~A�~D�T�#G��� bK��?.�8̎.`.�n��f��*��ws�Z�Pe��/������B�Ɋ���Ȭ�a�@��� ���� �c�s�-���|k�P_��{�2`Ӣ^����e��~�3U��������P��k�h���<=ͬ]0zxۭX���6�r�X�e��o|���m_�vt�Y|��)���V4t�Z�ŦP��q}yE�r�=�E}��N����R��l�,e,�@�������]O��-L#5��+"Ȃ���U���ryb�����_Gga{�%ۊ�h����>J	ǅP�o�-�Қ�Z�I��c�0�bC��I�p~�m���n-��4$^G��-pZ`���;%e�͇'��Y�F��Zf��T%�^V�:�6O�p]�_8g��e����[�aaA�6�(7���uO�����?�;7��`��L��Z��;)�e��!<��pz�ͤ[.��_���$3:�E� ���Q�
R�����!�MB�����_�*b���M(hP/�u��/FY/�N�{���~�!%�[Y�[L������8��Zg!Ę�`�u��i�+f�H���5�ju�]]��[��U��_�q�u�RS�W�_� � -ksF��Ū^�'��Ρ89T-�=�B������M*O���>�C�vܜs�bdT���z����2j/)>�
���IQq�ϡ�I���4�D�1wKsc� �֗��]�R���8j�e��(ѝ����Q�4s���ÄYFx����os|��_�h}�@-�m[�F�`1W�!�D��䈵��@�z���3!����!c��h��݂Q�2��8����F��_5B
�L�Z3��/����nk�Vy׀�eZm����6pz�K�?9�w�^**@��tUQ��JQ9 ��7�Dw6�cb���G�k�WElx��C6�`��?U{rm
Oh�y��^p4r��%��&��}ǙQv�s KҶ��VS�;cwf~&�����D��*�4��8�8���z�'��Ňfy>Vz���Re��Ɗ������s6,�
Ln��UCgɒ���t�oBv�[^x�=��'��o��Йb	M�|1�53ۤ����客�I�1u#XE�N 9�R�'#��-���9{"�\����q��u��r�5�Fc,�~�VZD�E��|ad
��!���鍁�J�j�Po#@�ʭ���!^wP�454����$B��wG��"���bWL�64��]�¦<��Y�B��dh�M:"� xb\�\�,_����N���ndtFn"�'���Yk�զ�����_��cV%j��=+s
_S����"�Y��U�k|0{\�y4�n������O}B�hBW�4��􍾖�R��G���h#m=*�@a�I|�m�']���"����������(Ԍ��r[��x�J.>�&c���E�/�_`>^�J4a$4z�oLߤSQ;�	UǑ�Q����E�!��ǚ���O��Qq�[i�NQto����Εxڎ7�Z��O�l���qE�C9��ʗ�ŏˀ%���x3l����/\��Q1����8���.y������N54[�m��q���xk��6����Cn%=�:z,���	_�4f'�!z{q���Ƈ��W(A3O��P�h��Q�I�u�9�u�zz��;_D~��?�����Dm��~��R8�k6��6@(o���P-;�[��B��&89ۆ�*�\퉝�j�h�R�,p������)����Hő��2̨3����L,Lm?R��6c�k5���lg����q�B��w[����|g��D�&]��Y�k�h��#P��B��e|��]a@�ב�~ s��@<���Mw����ڶ3Oe���9�2����q���ڼ�)���*���c�:Uhsh
@��,�TůM5OOC���zȿ�,��ew�`#9���v'H^uDah�d�<�%;l��Z����/�wk�S����T���=�K���@^�*��?0�����K7�Z�����]|���}�B>}s�8�K����h������z��E���Ii�s`.Nt��fl�mW��G*i��1!�j����]L �������1:��(Q��r�A|V %:R$T)�(�������)^�{�Дl4E��0'6dSzW̶�K^[���Gر��pH��30�b����+$tc��rKn�Q�\�-`
�u�x]`o.Z��w'���thzg5��1�Q�;x_�b���X���ꊫ\�>&&�/�>���>���	�Å�o',��"�������!��B���#�W��8�.�'ٷ���4����՗����.�O��_Nֱۓb �	�	�:'��煠��6����KQ�
!s�����6�Qn42kأ�� 2�N&��S"���"�-�$q��׆7{N����#˄��<�Y���>"��T����]���;�/N���?��Y��c1����	W,���ܓ�ϲ�PfIa)��#��?^+�~��>��;C��g������/��l^S���V�fܐn͔(�vx�iÓ���#D�'��֞a6+W"�%���'p���%" 1]�|�1�Ю�r4�-�^$~#[��|�C$�o};�)��[�JEE�	�����	��C��1���E�(E�Z/�������u�����/��k�_���..�P����^$�XԴ��]�������q�t�w�R&��ȉ���Uv�7�˹m��U!�{/.K<�uD<X���������DL��`s��S|e� zt�uzDZ[�]�T��.NT�XUp�U�8z�'(��~���J&�ʻ�ǈy��wGw�a����2�ET2	��3M����ƈ&2H�n����]���3a�A/̢?6�os�ZH�"�l`-J���k�����=�Ͳm��BA�E`�������#�ZǨd�N��>��_�4�t $Lz�J�n?{X@�����uup�U�p�i�(,���Sf�_�İ�����ZN�x�0�{�vdyU���~��~��aDl\�9}�|��뻪����t	��J������]#6�݅N�8�c}�N|q0�a��,1rQA��C��ЯY�<����N	⓿x����#S'o�� &�
��v��U����4�bN�����ˑn���rb`_�����ʓ�3I��D�����tF�HJ��9�%�B�iz'���ؔ�ðr
�&!��[�3 ����G"g(t�|����Xp�6�IB���3���"�p����x�/z��C�3	
��-�}I+�PG�Tձ��㏫��ǭ���}�c�l�����.�O�2�ۼ5��w�\o���}_�����X��6���Z�\�q��GD�6.��(H����_�}t	N�c}C�X�BƙPlK0��d�jdY���Js
A_�s�Nvh6�o���2j�  s^�c�t�{�"|O;V]��	���27� �g��*6����>���jO�.���#[>)M���	ď!0���7;X Č�ޙ~iBn��ؿ��Qzp�h���&O����KJJ��"(�<�������Y��pIr2n�)��]�T�݌��f�y�Yp?֨�a&�)��Pؐ}|,.�utk�K�w�$9W�a@yҀ��Ɛ��MQWΕf� �TK?h����֡�Gh�&����Z��1�2�>?����
��7������SSj0A��j�C'z������e�_�O��",&u��BC���.FVo��J<�	��m��s�3�\-ݒ7.����/,C����ٕ��������$����t����Z{�"�r[��\B�nG����{��Hg��\h�]G��}"�W�P�u,�Qb�;��d�> Y��ǩa�$z�uך�|�We(��?�t�{���<��y ����ـ�<��i�H�y�+M�Qmh����U�f<�E�ӽH��)Ć"�Ə#��D�y����e��S�u��De�Wu䞻YR�9����Q4.�8�~�4��ǌ'-�Hpd�UT���54^Hr��ǩZ��Ild:rNf��m2R%L�kF�7.z]}�ۥ�]��@��=<�1��+�Q�~��
o>�v>�@�M����|W~i9ں&��)���G%'�����%��zGM��a�&i,��y����!�["���4��C�2�'�i�Ԫ�,�A�7�C��q��*�̂<S��Yy�J�V�%����Ck0��yN��� ��%̓����&/��a̔)��x��Y�bUǭ2;D�f{���JF���{�p'�Z�
yW�Z��5ʺ��0�F���g��(=!?=dg�$f��8l�B�(�ɹL��I�V������<6ES��r3~�9h{�Mz�&�����G���˔<nٓ��_��0*�$�YӢ�Ã�P�`Q�j�E���S�o��ْ}�ܻ* p����g�\�Rz��~�>ضke��8p) /�I$�	Nߕ��d�h�>W��?KEL���Ḅ,ױU�t��o*�4٩8-l{*c�_W���s=�קԊ-�䭑͕
g��?�Z�y��2��ݸ��.���rvI	�S|ַ��K�c���7�q��Z�
��M(�?N��m��P59n�T����q��Z����Ù�7�3D�#9$ɗ��ڪ�헒֜���K���"�jp��棈V⸅6cjSq���yf�_H9��SP��`�Q��~Ũ�,g���,�jI=��a��G�'��]�K�xR���'��:$��I���8���9JɏJ)Ҩ��PJ_{Ԍ��&&�ϱ��V���>�$�+������k�O1��<B�Ǽ]>b�����J�m
�ي�(u:J��yt�v�=V����@���A�k��H}�}��S�
��ڷ%�<�(d2�q���ғ��0="'��MȨ�zS3g���e�%��U���2q�����\����xU����u�`�ZtpX�h�Vq�:�"�l��_z�u~	��l�l�c�X�Ĩ`�W�?���I��t%F�����`�D<,q1����ٮ$Jw�R�bC�_�X��1�n{��׿ܮ��$J�'Î���<���N�ߍpd#�Sˊ����>t�g�BH�ؤ+�h���m�e�v���
��iǟ;�8��S|�̈́��[ �t����*NKDut��W�v�>Qv6�q���6F���3����u}Gw9ݔ����;=G��L���L�|�W���N�]Ui��dM�MT�f+A�C/�~���-A҇ܠ��A���e;���2Q��|�?���$���L�g*<���53�$/뽽[�њ����Xz<�S��R�iB�1���0rx�M��:�]#Bٶ������!Pd�ܾ��9"��/��ޢ֏�F>����8���mpA@�߽36��Qba���n�X�3�Z��u=Jx}�ޅ�i>M��(��$B�Pj8����{�i�Q���BMy�y��7��=2v
Y=X�x���f���hol��<i���G�G�6%"|�3�-뇥T��B~c�c�ǥ.��-jW�O�ʊ�|�
g��yS���9�[���	��A`��C�uM"����������_e��
Nΐ7�GGcT����g����n۪�&�@��%ֲj�F�ֵڴ�&�Db��Ɏ�͗�:��DW�G�]���e�Z���t\���5"��t����\�o�m��$�����&yXe�t���\tr����`��3�J1�����7A�G�6��'�Y׎�>�%؟]!�6h����B�ь�0����wtN����iN��lk:H�=�ypĿ|��uy���w���> 8�5�]{�A#�H����Doi���`lv{ɪjbH�9��&��5��6%b����{"�I3�퍫>�7��+�(��g�s�a4_i@�*���Q�:�4���P��GO$n������@��gD�t����ۓ�r��i�� Ң���H�u
��%@�Q�|������xˏ��S�0�yX4 HU����cJ ۟o_?hW�E3�RګB2����<�X���Wo�^�n`��0����C-TڶB-*H�>��ɭ.��-���$�K�S)5�J���~��������<[�n���H�PS����I��o5c�����o�K;��L}/x�@���N�7(��4L7�2��KFGu�~� Jip@�Ťj�k�G¢��zt��8�W�Y`@�7����<�{�.V���k�U��"J����=GHl^��	#�6�^����<@���(�7��-�K�r3˺'tE���#�P��N�']���t�	�ۓe���"�Li�vݦ�Ǯ8o�ѕ�z9���ΐ�����{�eǲ%!��8*aՏ�Cײ��0�p~�!�2��|u�6x�R��ћ��/z���R9Y�>=7�$�xU۬�J����d��x��/�J���O9�ky
t�n��w^;�(��_�Bݿ�G��ik�[J�j���egj�o����j���O������[���nX��1�jG�
��d��˪�j� 4�j�e�ΥW�N�5*��k�9�}��>6��d��������-S)p%fR�ޏ$@��O����`#����W���z2�U�W�H)ہυ��6fw������{��$O�>�De���Av�����M_1l��QT�8��_&�}���PX|���!&�J���o.//�:U*�7�KB�"�jf�V��s�I)m�mS3>�j�N�$+'����z�f��o�ZuqL�J�-"T�ɤ�ɅQ�7�Ȉy�IH"y�3B�j��U ���$������H	��R����ݹX���M�|J��]�6.�)]�V� �� �|��>c��@T��ŗ�d3e{�R��Y)t*n[r#��o`.�[>kg"��H�ۯC�q���t`�$9����)922�ɰ�	C1�� ��� �tMC��M�[ڀ��qcJ�-��FE��"��Z��Y���>�M�h,f܆�[S��O�D�󋊩Q$v�w��޶`������L����#��ڶH���ru���ܡm��kČ��{	�TNQ�S��d��Xz��� jU�Ös�,T��pl?�Wؗ���ў|���,�8ї3���N�p���c�.�#������T\�~��6}I�=����;N���01���Y�]��B|�!�h	�����ߟ�h�Wi�����o�눶d��͈���(����F�:J5����&���=�;��0��H#�$�!��/*��v:�x$����{VN�A�ι�\n]�}���ǱT�ax�l�~����ɿk]B�\%I�*J�'SE\�;��V�RW���עD���E�AgQ8u,I�  �R��N@xj]-����\�#^�ZiXd -�Q�1--�\�9�NiU}�R�<�=��eZ� �xe�̞�WFmd�E��Y���Z�?���͵�rVw��+�7W�]�+w2)�Ls!��2��_�8�\6����L0��ަ�"�����?���A�*�W��Τ��
��k���Bm���nv���;��E>�(�(��N6�q�Fq�\#5?+�&��w|���c
�x�L�\W�<�@A]�]�(p���B́_�ۯ	�,��ᎈͳ&LT!.J
����|�{NC�}��qp��3�b�����Od�g=���Q�Ke�|q�ڮ.���`;������xtʔ"R���C/�#�!T�.����&A�Y����Hp����\%oq)(�NŎ
#�Ŀ[��xj�Sf�� ɖ��O����8�"�x�o�����'h�e�t���޸G���0��\
������`�����t���--�u�`7	��S�w,U���,�,R�ǖRɒ�ǝ>Vt���6m&*���{c���9v��6ۯ�:-Z#�rj4�(X��	j���[�Z���R�sU�'�(�.F����-m�q�GHu�8�d�ݙ:�����w7���},t۠�M�Y�l�ۍ	�]�i��$����z��V���M(F�N4��e����9�����߾$�*�5�/�#x�V�� G�bo�AV�9S���u���0����5Q�	��s���!�v�׾�t�a\}9����k���а����6`U�&�r��Ӂ��c��r��)�3�O�\�Bt������J�^�A>���}H������Ϣ`0x������r�'�y�lʤ�pl_]�����_���?]Z))�Yik�Tޫ�����*V��M����Ph�`�څ{�B3W��]9h3���������?�P0�_��������w|�Б3��=E)�p�W�@��B2�y�J�B)�?{��=ck�6��d�|�u-�6$8�o�I�
g�<���\7��qQ`� r��6%P+O�osf��=�ZC_aJ�}+*��D��������L��I��*%��=��\a����ջ�]���)�V:��u��m
(��߾��#1*/`����?�!H5���E���T�������ד��.k���i,�HW��cY�Be�lIe�v�bᚲ
ջ$��s��}&y~�
sbA)���^������%�S���'�>ش���lyKK����i��o����Y��b:�I$��Ic�7~Hj�u�cb�|�& O���M��9�7��b}\���P�/�l@vU��S�R("�xŐ&�������G���i��C�ζc"ڒ�2��tM�ؤT�����&��s��ِi��k�{�װ���z�$A�E�^�òr��N��3��|X�_�88O���7¶I�w�Th-@�#4ͷ.H��q5������N�t�BL&jIE�kc(9V�/��l���'�&��Ɖ������a�ZGi2�-��Km�Z�IF�NJ�-�;e�������HD�if��q����Y$���&>E���;؎<Tw�.���4ޔ�bpm_@}��5��aQ)>/��������SY\ǔ�6�����A�����~�Yn�uzX�3?��ЙAkD@t獞ƏV���!�=�X�����?��P��e�{l~kfkWD%�0sÈ������-����/��|$WF��z}��N�&�|\PXH�
����Я������1�"�y��dԦ���D�$N�����҂�'���t�5����̴��Bÿ��*���ZY��A<kSakrz�#�*bK��o<g��2v�{T@ Y���&���1��ݏ=����J$�9�?�D�&�)�;�N��!���y�a�y���bZyǔV�Z�k�2b��^��o��3\����z�Q���S�i�k��K>�__�a�>~��mD!�є�p	��Vq��<;G��q���\z�ϲI6Q*�?�� �RF��)�Ӑ��+���O�D�M܏��ed�Jԁ��D
�7�g�O�Bd�5{\�V��_�`R� �T��"�\WA���F��{�f�<E���qghK'"V?v�.�vz�6*�Bz\��a�u^d@�A�r�?գ��؜��)-��v�C�\�h[^}I��:��~���y�c��2��|�������W�hT�љ��~��i�zTx5�*U�0����r��iT�!����B.����8q"��
y�i�"��u��/��|M?�����m�^{�>���%5�z�~̗>�G��V��ՠ���[`�\RBÑ����˞�a�(�-�9/�  &�����V�������,����Ԍ~�+`�a���[N6���5rTT���[n�(����a&j*9��Ws�:V&��F�'4?´�?h�Mѡ�H�Q*����)�SԹ+��qN-�Q��<��Fjc'0�Z�f�v}\2~�G�[Kx�Q8������,e��gÄ���1z�՘��[�oO_��y��*t�#(z� �2�힌��y�f���D�f��~!^\qy�D_�ks6��������2��"�g�p�G���
�y ��IId�)|;9��y2��ҳ^ӭ���R2�񷾭S���Ӈ�f���I�d��P x��kuU�%�&Wʜ��V��5���Q�	��i����`'O���..�0�����L��+f��#D��`t�E�*m>���"����wt��L��:"p���x��n����)�f��Ik��zئ��_�_K��z�l� K��'����^�
n�N���KP
/Wn���xyHWE�����qT�Mm��"vV��e��Zs� �޹-���tB�{ʇ����]��r����ǯ��w{�|�vG�[+�n��^N�O�8�<����|�#N#�8�n]e�S+�o��b���ڪ�D�p$�^_�\��|��J)�	�-mI�@E�]�{�?�s$msң(A��T��Z�K{��p&�9]T���e	WĮ�1V�s�Ĭ]Za��@>hl�X�8I�kRl|<�j��l�z�"3>>~d�m�n:X#H�Y���bE2J��u0^���G�r���d�0���2��y����ancW1���/J��"׬�8ƀy���	������wr�/T���ݜ,�H�µ��Ƈ�����/��U.�<_�}(�{�n�uv1��V�����CF�4���~�b�549���7p�s� L�l����GQ�tP�V��Ǯ�0�X�߶^V[
v���Gak�K0m�/]:�z!f&��;��7ƒ>ޣ�55��3��<}eT���Ipwwwwwww	n�]B���;���!���ep��8����߳z��]�w��!cԆ������������N�m�F�Fξ�d�j��%8�DHZ6~�B![�r3I#��kY���)��ߡ�P�<�3��}!��e�D�xqЍ8��<�9wpP�	�����ߣ����E�}��6g�Z�X��S��ٗ8����כ�aeUS	�Q%�.���	������R���a�y֙0�����(�wB��44tʴ�O�,�\_���F]����'��� �ɚ�����!d3����]�B�e�p��]Ґw?�jAG�bW�"'W����P*�!�wE���INOy|K�����G<L�4
�8枡�(S�n���������Q�����"�ۿ}��X]W ��\���W/�Ds���Џ�@��J0Y��9�	���oY�]��'I��s��u٘XZ�e5��~�|;��������M���'̿M�C�R�X�^�K�(`��g(�w�x��"��g���WϜ\�/CU����3A����:����]�3˭����������B���`�?��,<��O�p��Ǎ��S��C�4 )����b�l�W��)�3n
��5����J����6�',�M�J��ό ���_B{h�8q9>�����v�fw�x\I	��7q�[��9�����7��v�X6�� 4_Z����hY��ā:ڬIv>�a�{���Y��6���Ne����U�0*���d��?Yw�:?xi���R��t����I�f���Gbx�[ 
�)�U��W�����Q����Y��H{�B��z�f�|L(BK�)`C�D_n�����9]ߒY�5���9n�w�� ������]��Iz0��L�� �BKjr�	�G���;����+�L$�bg�� �ko�Y��:��v]`X�m�+Y�V�5���R�����#�l�C��5��=.��s���ke����z�;(
��1��`�f���(��m�y!�d��	�F��
�2�v]m�:����L�)�������/aq<��9�܀\��?/k�_�+��c�M~r�'���u�LYd��k�C�Ҋ�cq�6�������O�bMXj�#��c��s���.�w��5�x^��e�U��a4��ȳF�^�i�\k�4^Nv��a�?i>b�N��^p��No݇45[���+ #�C�3�^��G���\��dF䆏�^W(Q�I�5YR�,QlH�(���<�qh�b�N��cR�@i00\�׵�W��{�?c=Q�2)��t�����M�I	�P"S��'��N�2F��[5�;��~Œ�x}�|:�p��}l�c5io$tF�F�諺�j�~;���K�hoc�������pf:	���j6%���)�E��ſ�suUMr	
���"'����ƶj�T{���dzW4�y]��z.����V}/v�\�e,��㗧��),�c�X���S�=D�����v���q'`��p���k�\A�5_ˮe�������z�-{��m���RZ0�_�^VN��ʭI�e%�	�K���tC�8a�J#U�J���$ky}��u�����*�l"d���-P�"��9�nW�,�G)B�>�~{��|u�K���,}c㽹r�
�����x��?�p�'�j(��i&�۬�����)*
��*�k�����m��WV���D��Ъq ��\�-��A<��[4}�;�ߙ0��~��q����FǠb��������ګ1����^#SCMY{����B	�"�2����|�_)|�?��a(�%��'��|�?S�.���$��ϔP��21i��v�RrRrZ����r��	�(999O��r��'�'���6�w-<�{�;]�c%o^����Z��h�z�y3�Z�|���	�%{��o{d�X�p2Ș�լ�5�^iyXy��L{��|ߦ�*�H���/���w"��Ȓ�,��u������C�:�)�Է����я'�wuIf�쏆h��TLu����r�,��H_��o��Y8�~Mi�8!�\#��x��Z��9Ec��n'�xH�Z�,c7_&7wZ�O�>--��l�0�=�ߟ7�UF�55��T�� �z����G5+��<5��Z�T���ԑ�}S�y6��u|�5��T�F�m�o���X ���U�V#x��4s����ώ�8V6&r�D�(�����앣繣gܱ����Xt��}��!$��������gr~v�>�UL�H�EN�z�96�8?��3��!ih�|�s�&{} 	�]es����i����t�}�����m�AVJ��_�Gh��9��5v��)���`_�z���	*��B��&U��Ll9�F#l,,�PC�F�g}�W%��rL�$<� 㸖�������q��a��]�(v�i��6qZ��i�6{q�.N�KH/Y����{�K�#ϙ�ڻ��B�xR�l\"����ވ�[�׋ޠ1`]�/�4����܅b>l��dAfdL�B/b�s�-j�ɖ����`}�Hce��̘��m d?�����ǯ��0r'�%)��`�GV�w)���̝���ɴw��e���5�i����a|���g�����_9b���㯸�J�zc��<NM��?w��ʥ{�a��r�T0�Ybշ�)�\,<���}O�r�C�BB��N�˶yuuu������n�'� 999��b��!���A�k3�#n|߾ƁY^o:c
D-v�(�"�1J�t�ɺ�ttN/.��7;�[6pe4���6.^N^��g�G;�6w�z��L$����ܛW�ua
~ ��,A+c��B���o�b�1�̗LL��OLW�u��x� ����I�S5[e��7߱"V����W1ppĺ\��g:6u����U?q�,#n����Vݿ��� �9k�bf%���<���r�,k���S��t��L�Pt�E��=�8�hi�]Q;f�|�kX��9o����������*5麁ѯw�a�Z�b0�@�s>��/,WT��:i!�M��6ee��S#���ּ9iZC�]��p�`fb�
>�A�h���U��LH`Gd~��3�R<nD��/+ܮ�咽�
���S�П��ntq��X�.�py��a796�b���R��]lk�Ri��C���z��+0�>֡\H//��D4�q�1�6_lJI�5����NG�W3�_E��&0�H���%h��絥�Q]=�;=���h��;�#�K���Ѩ�H���dD����UO���^�S¡b���7�Λ�ի�������i�\��L� Q��8��`���7��Z�vb`m~�gޝz�j���cԞ�'�{X��*y8mPqO3F�Kė��&��mz 䀦:n:)C�ƹ%�M�[�������r[Av�wL@x?e{�N�����k���w�v_>�n`����$e��U�$Kt⤆���whNȸ�#^}-_ %��b_�Dl��Qӗ�Q��`�	se}��e�;�����B3�f�(��S� u._��J��¸4y���p�R�E1~2?�KG�x.x�;(k�y]�J3�y�q����4�VG�G6���V[�����VB����l ����ZV���??Ζ�DON��`
Z�j��⃯���:z$D��|�n�_��G�vî���`�'�Z�qy���׻%RF��v�#�K�S�3B,"{+��%�����S�'���ZI������5���a�*����>��kg-�����ou�M��=��?����]����y�s<��v�+�z]>�EV��lf%s����M�l���(-�?7O���ls	��8=;-𒖊��	�oEЦ����=�]O-���Ռq�c�ퟪU�n�̻�D������"}�c�	>n��^�����,���R�]�?���I�

�D;C���)��?�;P��$��O�ě��e�#�!'��j�PVC��"�o���Wے���,�;K	���;Hw>�K�!�*zS.|B���Z�۾�[}�Hٲ�.WG��,M��8d�Oŧ��x[���{��;�s�D.'k���p�˰�W`���+a��V�����FMm}�*�n���s"
���%�n���`�׫�=̴��2�VD�6�:��~�ivѡ倫he�VG�Ac`�u:r��W��MeTg�k>,`}f`u��lyd���9A!cM�R���6��4h!È//ƭ�~Wأ51��ōc˾~=�x?W=�g��0����>��c1��k\S���q�yZk����E�EO)����t�_��"�'�]<��"��i3��ʱ!�4�%��e���O^�?�] ����v}�"�q����<�ܔ�Z�������FDp���ba{�~�xg�b���5���g`���q�B�~[gNѴ�SD|�0�)�1�Y�&i�^;�c��C�4�/F�y[(���妾���a�EȜ�(^�������=E�mxW��C;�����
a�r%V� ??���Z����DmCA��@$!��q*�1A<�f�#v���[$�����������S�7F��r��_	�PƩQ^ʼ�h�d�]�+��7��@)�Q����ѷO?[���)�����W������6+��r2�^�:f������+4����\l���Y�s�֡P��~���8V�89;sf)gL�T"�Է��:���AO�Pg�+��#ە%Lqde2c���9�|�1�P��R�;_�����r��b�7g���X�d�G�����Sv58��o���mˠ��G�w�b�=���m ���?�o30��^l �FC����#B�tQ�?LL�>HX�#���lqD�r���a}u��A5��T�V$�(��˨Z���m��f���?�����ͅ��$r�X�̉L=�F&�z��BZ��_9���vTX(U�&�Y�4Y1�iv����`k��2:����Dg��0�@GJ��V��S�M�"/r��{�{��؊�D��ܿ� t�α���L���t��:��G���`th�U0�I�2��Obb��ւ����A�3-X�(�`k{ś�oZ�X�B��-��KeB���P��;�����a#u�"�����v��3�8wq��O��Zf$""��G���X�~�=��SZ{�!�2��)Ge�0����CY th�x�y���1O�hPu�*�ut.�S��;ډ�+2�E��U��r馾
z�l��z)�=��4�ߝ|p	<w�A�%�b)"��k��?��w\v��� e���5�y\q�왮y�9���||�sX`�S�&Ҳ��r̸��r���r����\���u9vR��/`�2awB�kC|~U[畲M��m�sP��"0����(+���>I��i�q���B�Q�|�����Z�� �&2�G�-ӯb�cF`�.p�M'F�X��r�e�WV���|�"=���z��3�#��\������Ȍ�btfs_Z����紐w6il��[=���WUYʉ�*ҝT�V�z�1�u==SN��`b��^�l2(��:�����2�VP2ɡ�p���]}�i��疦���O>K+�gu�R.�5�_d�>r���2�x�%7��:g�5ڦ��	�ok���1A�������FN�$�j��E,���B?��g !�oͿd�Sf�q�=F�A��t��TA|��������mM��|�nh�X�_}�,}X��R��S[eiyY�AG>L��.�WI������CE{�����������t�%�}�� QP󄑽�8�$�\3}J�?��	C)6((����`���B&��3���!5��J�Λ�o�oI��f�nP}��p��î�8i8���S��2��[oA,[�Q�Ƥ�;t|�/�@��"q��N?�K�u\�k�umK�J�ࡒ�ǃ����q�����4�w���������LJ���Ԟ7x5���_�Q�;Ee�/�D����Q�ñ�m�����+��[3_A4g�̦t�!��Ǎ�^?����=����T�o�L3�Ka�����Y:�hp��V-��V<���Է��-�B�oc�O餪d~�q\o�o�ۅ�$Z�g9_�{K �c�C��)��d�boݐ�����3�{�ފ����U�o��*�j� �K��`���y�^�<T��V��)�)��N�x�C�����jI+h�Z����*8P	�a�]�&�e�C{��o��[[�;�ҳv�piޔ=C�,v�D���<��2eu^C�Ҏms�������:1F��oK��<a�e�W��;[7�,�[����@VA�^�fZ�; �P��`P`��7fH4s�`7ڙ���P[_��j�	�7_��Yː��@(�;Қ���G�y8	�����̖���U6{���Ĩ�+�c�|�V����r�]*�-����1#��l!�hz����L����{�X4}��^��3����F�q��p4���|��.�|���n�.������H������0WGeSldX���J��8
!�@�g�Zd*��%���[���qJw�������� ����!�1`M%�;����p��p�	�7�&�$�$'Be |� �Q�[�T�b'�*XB0_�A�2#��e6s�R���4+Ӣ8*���i)���1��K(��;&=�׾S#6<�3�M�\b�������u��� �����S�E�NP>b�ş���1�������vAi)�d������m��8Y��ō @��ZOW_g[�]�� Ɯ3cb�͒*\iNV��s?R�2>���;�츣$�9�Na0�a�
@F6�����,�yw��3�q�Ԭ_/R�Z�D@�hq<�W·$l�i�{��S��Loo��AR�2?���&Y��%�Ɣ��s�1���ODU�n�4|��Ӭ�>�I�T���QYSU��!
*��J+����rY�	.櫹�x�{��b�.ƫ�9fU�m����z&A��W�y[��ݪC�8D�d��츙[KX�Di#"���$MT��l9I=\]����r���#}��)�����F�p)vf~��<ɸM� :�؆���Ee5�T
�rISiʻ?^�p@��w��썠�hX~/�K�qR�R�d��%��V���4q��&��9��p;�;&&b��=_��t�<4�mf�酜�����ɔ�޶B"�ѳ�Mlu�������������0i�� V�C�$J����}nMdNg�?�i5��o�h骒@=lz�����T���9��_����W��{�����|�}�_�H��0~p���*�7W���@��*��8�99����*��-
�q"�#�5��$�G���U�LZ�Ά�
���(�b��7	�"{��{���0�yZM��
��(��[���=O����WKEԤ��L�Ә���V����OnG�'�3fл�!ؐ��Ԟ��n�v�J��аE�g��7I���x�����oyN=�3�p
\	�9�WB�i�Paz@~IlK>ɾT}���;"iD����/)�|��~ER���#� �a�X�~Ј���ېn��R������rd!WH�k�ߛ*�������`�.�&�������6���Cz8d�X6�"�ߣ����9	�ʾM�ķ��"�u���Mƺ���>Wpn�F���o��v����R"^��_+U�zRZݍڵ/�i�9}��$��dM�j��M0�^�8�5���Z���/��ʣ�*@(Q?��&��<� ��ֵ@[g~��%x�%�'��˱9�B=�5l-u?���%�h�:�C�9����������N ��|h0i$�d�>��27�0��v�J������w5�'#��cE�J'����ؽ�Q���fY�&�Dg�O9X�dh(��fa���h�tfx��U�K�Y�; q����M��_�$RH��J�kDs�wU�p�ճh`g�Wo#�0�����D�v�l�z�[��������^�+�mk��n=u�ӂ��8Q�*���a�����Y
�pf���b&�.�����"���_8�Y�d�Ӱ"|�u�����q�V��!գ`�tnf�p�0,��Z@3nE�2��go�YL#o��W�|78J/`�8oV��zuW*�|Y=i<)o�ꛐ�i/�=�
���-�x���	5�4Ƨ��y�F3 ��ڻtux,y�̭y���j?4`�;0��ؗ�щ̃�Y`���P �8����T��ຣ�������R5*���"�%��Iխ��RD�QJ���3��`E5`�J�I`q�p�٠Cs�U2g#���z���H�,�M|�J�>p<A,ޗ��ewS�W�')�]�]���F<�(�<�Y�|������p�gpy�>s�ׯԛ����~���$3���Pw��=̀��X~�����x}�B35f8���C��^��s�i��9��!��~1RX�@0�Uw!b�j����w���� �c�@���fZٛé����%�;;��'5�w���-�!��Qt�]��S����T��=E���h|l$�j-�1Mid�l鱨�w�l�� !P��c	����&�� ��E~F��2�FrYvi�t9�j�hc#��qV^�~}2 ��g��zh@��Ή UdF�{�d�Zv�a��pH�昌3�ĒT`�o_Z�ưP�cH$08H�0C�0�u���Q�OĀ��O��Z������8�E��E�#£z,Ěh��ϕ�������5�9�E��|���̒/gL儮�q�b�&<#���9:*_xq�VBY�cC4-*�h��i�pO�]����wv�ה���4W�ϴ�ymߣ�S1֥���9b���v z%qv�IN��M.>4\�#_w�ߑ}U;+�Jx9¢���ӻ���(GDh)��m?��Ӱs�X]�:�����o%!�y���$��/䜹	Z��q�yѤ��e�!�_\H1s:2�دX�7S��bN�+7YнaD��ᣓ^(�@��% PK�i������$�q{��P�y��k�µ�t�:�$���]e��"�}eپ=�%��[��#f���B�&�Q�B4D	ӆ�Ї}ٺ�n�5�M�;��e���k"|��wj��@6��F�v��r d3��"�:���m<I����r��Ӌ�i	�Z[s��Ԗr�J_5I�sq�!�'�T�%���6���K�8�RY�X����DE<�������rXw�5�;�IP��p��*ˠaiZZ��z82�Z �K�B[�D8�S��x�GԎ�k�{�#����
n��ۋ 0�M8SFF�Y:k��bVO1�_+��o8�����'k��յl>�Қ�-;����	>r��|�����2r]��%Wv(�����ˤ�R<8��J�(l��N�����~M�x4:��,�'k�#�<9_	����:D�Tn��ޚ^���-�O9
ʞR6��j���}���MX|]յyZ��%v�	i�,��4Ewz��!�Z�Og����J����V�����.��L�ϖ������\�{!�9������C�#�᫬�F���������W�|M�:�_��=�U��1��1���7�[�W��K���D�E&Z�X�;��
�q�٪��m}��_�[�/����|i5���no���N�I]�s�9�e]	Kd�2�}�DF�+�ƍb��#s�ǉ�����rhe�qΌ�V`�(���ϛo8�BQ�;��f���? 4�&�K�+i�~����������I:��j�l[�sɰf~Q�R}��l�nP���2Ti��TSJ��<N����_�x��)�VS�p�:RL�W<,O��m��ۥQU�}<��%� R��,�#��Q0�Ft��bۄq�dI���p�f\�j�Q0GT�gi�=��3-ѽ�1������ط����$G�
���{����#żF9�_l"�������$����~a�#:�(��T�T��[�[�Lp���ۮ#)�z' 5����'��xY��t��\�t���u[�,3�:yxQ�ZO���HsB�(m��̔t���Dk�Rf�+���x���%�If�Y�@�8ʃZ���}ȩ�T���ҙ_�E�o�`�YH��Q�8��kf�%���oNN��c墕���[Y��dC;��n��20N��`���͋쾙��\�	��.X��U5z��Q�5=cs������њ7k;����G��<���|�	�����x��<�õ b�RQɂ���Nؽ�a��@���B�ʛsSd�S@�hu�ޢ��K����G�"����֡k�7ȋV�bL� 'A��*S���!�{�-��?��l ����uB�h����l��|���Y�5�E�-���O�!T�.(�U�7&�������<X�S��q*�}�g��hq�����I߯5T0.6~B2lf���r�4� e� �
4�I��By^�l�u�ם�R�1a/׊�GO������r6�GE	j��2�����F`���ph������(MY���goo�χ|���?J�Ы�Q�I�0��yl8����.�v��5��,N<���G����do�+B=��OɊ���ɡ�JCш�'޿����k������;�Y(��7e�.niE�9	�N��\��6��$�!0Vo�W6f�/-����9V�vT�����r��,�	Ux���l���dSԹ����"j�������x�j��0tEN���B�X9˗i�����!�OR�c9�(%O��:|7�(2��H����4��}�/A��ڔ9,�jd*6O���o��eEWq[�o��\��v�Q��BX��!��-	���srf��V�@�m0��L�'��Eϱ�\�}�����<=#|<�JS���~~��3{�{G�OIًo�YJ�]�̚�O���>�����F���9��**�����PQ��c��m����y��q:���#�$� ���	[
�7����w�eLq�SvB�:�Ƙ*kj�r�w�	�h�Up�tt�"�{Ĝ�Cs./AJ��V�e�3X��W�Q[~�R���l�� ϣ¼�荗�Z�@�����N�5L%o�u��;���!v�P끬g��R�τ��2z�9���o��������v�Zӈ{� `�1&�!�N]!%o����z��<��znpjL���g��G�@I\"74?+�EU|��&����NX	����$�U�{�2��*��.7�p2�s["�>��P��9�n�D�������e@`�w���nI�fC��OR��d��JE|~e����uUD�a�����JM
k��A�%�O���+�+��ptt [�PΛ���f��4���9k;Ң�o�u	Ѳ#�t3�a��	�~�_04�����n��I������U�������4��8�ͲG"���i9x�r��S�ˁfxM�é��w�=U�V ;��I���x��Z�Y��X�`7��C�����h���5tJ�r�Q�L�,���N8���t:���V.>ʕ-��;?	<4�ll?!�����g�>�D�f)N���h�Ù���������D���8��
}�5��H�4:Q�����[F֤d
W�ח���",�s�h��ԣ��A�R�l��9X�>�F
�g��_�3�[`d6�項b��Y+)��)MȢVV@]5؟�>;�̄e!d�!�;�0_�y�m�������� b�˕Z��&
-��U��?'D �A�t����l�C�Qؖo'$��	��)�`XX�B�mh��pO>'���?Y%��k�Hf�� 7�'+B�����0漅�%3��%��ǧ��M�_{��D�)��q.��c;p)���I\��r�n�n:�V�vbr��6QsO>��`����ƀ��.x �|���~-����`���n���^I��6�2��m�Q��� X�l�y�'�g�B�i�1*�+�?��Z��hv�]�)�� :����p�p� �����O�7��Ʌ+g�~�>�"{�+�C����_8��0je��Q��8��I�ZiZ�Q���^>+2��=�g 4*��8s`H*�;}c�x�&x3����ԥ���*�y�@aW�"n6��J�P�B�ۛ���X	�u��������ɸk���-_
�ʾ.�*5�~,���}������9�zk���`��ڸ'� .YȲ��W%}�<�N��T<%}7�MR�HV��W,=W	��o ��7=�1Ђ7��V���5��h�\���Fn|���0=X#H#��lhҞ�4�O*������PA6\���9/���;�;~2D�e�y�����}�����N��X�t}6Pѡ�KGc��h.מ�Mn�2��(Z:���%�8D�(�GvS�7��e�̒�@�b��ph�������ꨔ��+�Ii���&�=�l��nU�	��3h�p���".'��8�OS�w��z�<J�6��K]ֻ=",���K�Ԁ~�^>��5��BdV�I}�|�L%N�X�X�w�$�tL AR������4aY	g^¾�&�֠@�4�oB�I�	}�X��-��mල�������M�s���I<���&l��e�F�5\O'�@�����$2)������Cąϧ"����Otd�3�_���q=qҨ�Eiq&ےRNJ�����c�K�����X�tYl���[��D� o#֊��8ݫ�6��� n$�w[�4�� ,nI����$D�|��**�B� tyun���O����>=�����.���z�"U�2R��R
���*QՐ�����]�����|�GW�J	���Y4om};rZy p�ۆ���%i�����I5Fc�~'�{�6��f����+4z�iA�i�C��_�n�!���/�w_�N:�;��]6Z[�U)R�� ���44���C�{��7�*����W�3��'A��¨�i����Q����6R��l[���{�1OA몥��W�\�B1�?���Fqղ��g�j��L=������Nq(Yd���(I�MP��I��땦e��*0��,����ËƖឧ����&��+�P'��&�OV1����27rғ���瘜���	繜?y&�援I<��Db��g^��Vc�!���oAa��&�OZߦ�މ/ܱ��<'z+���&i���
��7VG`e�Z�s�/�^����~��'*�pBHl��n�V*�#�u����k@�wy�|���u�j���yHܮ�T/��7Ĕ�|���D��_�^Φ��ٲ�z>�̵(���m�f��ٰb���/�F��MD��K�Y��/����F4���W�)��g�U���x⣡E��K���F۽�0��-(�<�=Q�|+�y��Ť_,�,o]���R�������U�9��4�+�g4�0�U3�n�����8.ʤ��ߦ˄�Sl<co�"x��Kl���-��-�t��m�L�z�lA^W����-}0?��톡�a>�u�΋�m��
��j9I��6��C��EV���!u]��&:Qb*��T�쏁@�]���b�@�6<�qn���ۋzf���ȵ� ^��x���x8�Q�"QS��F<��l8�.T��JIM&ʗo,cՠQ�D G�}R�0���mbů��T���T��W.�pO��+|*i�r�b�ԕ��i�MZ��^ʤ��it-�\W�����(=�O�J��Z7�9�6�-v6CN�J�*����",���!QQNd�g�͎�<>���r|2�蒋��������nʚ����Q�fk�]��_�m{�V���7v����JKH�>8�Rd��	m�($����5?�(�>���ia���>���1V����q>TD_ t��,��H�K��n-Y��7��rM�g�bZZ^��9��D�r�gU�jj�N1��F��	[�G������8i�c:T]Q5� |,�����X*��í��V6	�)))��lU�\��4i,����	�M�Jў}�3iő�ӵ������@�G����Fi��ee<��/��i6D���ic�pPx�����U�%��#$I[�1\A����O��Q@0#<������#�j��U:�-A��+&-��д��d�g�������0s��m���u��T\}�`/��t�6��#��Ù�Ueo�S��{�Qf�9�FC7.G4`�8A�.d+��3��P�Ry��ES׫�j�"y��
�O������(��蠟�H�� ���eMdS��6���ȓ���['�豑�x:<�'�J�i-��WPN?H�M�u�G.�#4�bd�M����ґ���2�����\��C��� X�T��h׉Ӏ,E�9��Ԣ�@^�=�p4!U��b���m��w��P�&��/>{x�!��;ADȲS~#�fAZ�
sc��֎mb�x`�8t�睬�مyd
��(n��I�����	�a�0�&9P�@B}�b��Z����C��w|&'Zݭ��],h���0+}�f�b�T�d�Q'A)�DP��Q!�ʞaJn���[/k���L61�h�,��#�pG���"`>㤚�E�ti��|�]����|�j6��|�\�z�^Rj2*� ��J՞r�ѵ�@
���H�V�)h�G(@��qO�-;����~�r+�u��<xN"?�xjhKm�80%ɇ��S��m/:AR�s^��I�%��ɫ~D�Dn�ʏ��B2p2�F�n{4��E猡��'prq�t�)����8IO�<����4^n���hGW��b�^��5����b���Zs�V�3<�C�7��j�	2N�rX}v�a�`h�9?�f��}K�
Ӄ�A<�ۥ��鳓Ņ���U�L�;�r$^����"�E�ΥP�Qm���x�M��W�x��싈A�f��A�O� ��k9��~�02��I��^�2YX ��9*j�G���m�g4��"�Ҹ	����	ڴ�)2%� p��/dP��r�Li�	N�cl���Oۉ5P���n��_�\i�x8�,G~GA�k?<p��!�QC�>=��
5VoӸRGI�V�Kg<���jM�'[G�Y�אl��sZ����ffR�:�Vj�>���ͨ���x��y�bח
��H�
���uM��_����&cvb����O�%U��9>������Z;�wTZ�>��-p��D��v��Hu�J����K(3�s�E�Bm	�x
��>�/~�t��&�!�/w�4�#_|�����5j�H�����͓�"o_I����4o/BNȃ�5��!��:FR�K	�2�i1]w�� �h�e[6��:�Rz�d\˧���g򀧋��%+��#��R�Z&�ҽ��EL{��dߋF�Ad.���L��_�'�Y�� U�f�z�Z���]���bDGZ� ��Fp�䘝t� �Tڨ.�r�k9
�C�t�g��cʢ�G�{gN�TZ�h�f��)W�9��%7��6���j�hW�v��0tq�W���'XU2����%B��Y���&Z|�*�f��u�Ms?�c���ز�ZU�9=��Q��z�/�w��(��`H=<�����20�H<w���t+��QE0��9���G��xp //�m�c��H�|v|T��v�g�
�!�`b6��K��I�1�&���m#U^������W?s��ܱ8?�����s�^����S�4��\��е�Kk�nɝ��[n�v��D>F�@tx̢�����p?$��`���A9rx��n�g���? ���(%18��u�C�Ur�|̠A���Ƚ�c�/Iv$��ef(��J���hb�.5�b�_X�4����Ơ���D�5��=ҢwH�J�@C!�	G!]p��@�_ ,�@�Iq���7�.�K�����W*	�|��������7�N�m
<�o�h��U�/��R>�Fd5��_U��v_~�=;����K�qzqAWM�����OO:/�X����"���*��
����zY�yG�pdJ�O^��H�m`C<D7���:�{�������#1P����L�$O"�u�g����峹1�#�xvRC�E��$j-4��#ݸ1�EM�[�ѳ��*=��]~��oA&Il�ibZ��L�{�z
�d�y"'A�uXq�dV�5�$�g`΀/�n�4ad�w��<�G� ?���|N i��(��!�Wy�յ�o��i=���:�d��rnX��mJ�S�[��Ǡ�%i&7$WT*�(�R�K�����XK���0O2�9��q$׹�����u$�:Cu��'�_�{^�Onʑ��HnjuO��y���?ؽ�8ś͝z��˓<�Aش<��;�Gb,�B�PC,,+�C4;N�ctL�6���������!�>.�s&�"Th��J��H���B��G'��D�;/S�C�����1Wʇw���`�[C� �#L :�Z��]�����gRHY����mɟ�ml�7��g��XS'��"uN�M��Ai٭��T�����F�s�o�4z�D��_��oB���؎����k���t>�9r4���˞�y��<�x�N��Yc�?�@+ap���?�Q�'Jɲ�G�W�EՆ[� ��0RCwwJw��tw��CwI��%�9"%9��C7��{�s�k�{�|�u�g�;>$�px1�'P���Ƀ��𧧲c'��j̨jTd�`x����@�I�����7��Wm�9ը� 3)I)���8�Jl2�NH�T��%p�S߼���QR�}��nL��,5�ɢ6�؎ �(��,S�2��}��*ptT5I�y�@O�(���2��}��~���ѓd��N	���$p!�� Rt�g�$UCL����q"��l�����57sv�ms��뭹��؇���s&�8v�p�\�IT�H%N�wdtG�v�E�Ԓ_���Yq9Ŷ6BN��3N�s�,�,���2��V��\؅݂��Ņ�)�D3|y�Ej�܎Uo?��oԗiܤO�Lt��h]+��X�ƭA�I�֢0�o�|�B~\�Ku8.����L$���î�Z'@�\�"(���҄��ܻ2�N��$�-l�q+���.�#�լޥZQF�<:�
A1��a2#=#\���ǆ�14���M�Pnn�Jg��$�>v�h�r�{j$�D���j���r�%�A3��9S�fS���k�MZ)�7\�UD	z�"}D���\sKCy-9�+�Fߡ�e�<�cq��0E��K��a[��La�(�j�zJ�UaH��ys�wa&P����"f[��X��x7���j�\�7A��� ���i0Sh��|JO���h�Eҍ0�p��y¶���}��u��3q
J��c�ư��&��K(�J�������k��(��a�ј���e���8Q�Aꁏ�h��N�I�c㱠n[�G?uϴ�p����.z)��5�z®��������u3�6�+�~ʜhŜ�|It<��7(1����Y���2Է�w�Sg�]S排jx�r�uN\\�������Y�I;}cv?׺��	�6~v
��q9q�DF��=�g�Ź�7���x�(q��,a�z^On���P˛�����H�|X`A�!���K�Zq���n�~�����J~F0���`���0�P����{�ޞ�v"P�v��۹����9�T"�h�{��5�B�)&��;�Ӳ��}�c���H�X-VS���v�tmE��t�y�:�@��PU�!���\ ��x5c��7��a_�|�&flb�p�Σ��k�����α֨�h�g	�&<%3�ٰ4M�3l��g|u|Bȑ�!�~�G4i�H�Ɉ�����%��>�i�1՘M�#>�dg��ꂳ�A%6�64�p��O�kl���9�?�����+���dΚ��K�i"3"���s`�-����KF~So��_6܃:Q�E�x��U�,�rW�9��.�T��V��3I�}�祈�a��ǲ����Zr�K����=��RD��ܩ�@F`�j;�io���)��R��zO�b��/N,��a���/��.����=�0�Ҷ]�
�F��(�izN����D#�l!��qO�\���;���"�,���(�a�}m�����E� Ub�+�!25�פ@f���QIg#S�7��af�H�?˚��M�����TqWVv�si%�+��V�<j�QV�u�1��P*2�ބ/��������DbYd~A�AR3ݺy&�JFa#zJ��L�28/�h��&���~�	#���G�K-�y��a���S�@՝i�r!����g��Y�H�S��p��!�$cei t�V��H���D��%��^9�B��BK@0a����E��~7oo� A��
����p�ap7NW@��ýv_�	�ؓ��{5����#����T�(�������I��s�������؉�]q�,4�!�UP��l	������߹1��P��]H-� �2EWR�=g��I���>ڤ'�@��c����7%%�*���Z��_c60�]~��5��:33�26OhO}�|
h�F�)�)�A#��$觘����2�/���׋���62�e�a�^�m�W��b���яl�qp	l��(�1\�v�7]�3�d7C����w���A�U�o'{��i�..�5^�u��
��p�
fU��	
��;_v`�O,�0��۬����>s�k��}]�+�C=u������<eկ*��mY�z�>P�aHӛ���?K��0Z�E�I��꯷�m�C�d���a��;�\���QΟ��iұR3[O�o��>8����Wv��ԗK��PKJ��}Xy[�c��|�J>>��������%����[�}܂�/ξ�򋊊��T3L�N�Z�j��7��Ĭ��_@�L�f�^%������ {��6k?�Y;�v5��� 6B�y��Xt�[#�2�/U*O=+��ۏo�>>�.�o�?d�-�@�{�=o'�c�&�F��Q�&�����$Ľ�K��|O��k/�`G���n��F�iC�m��.�3g������ �󕚋ygC�bW.א��)��N������9���+")��$K:I2�޻��[lqKOV�0����L�<p�;hƓ�`_���Dނ�L����/|�_;��8����w�~cZ�q�= c��<��<��y�7���3ݞ�Q�9B�I�*XԞ�jǭB��v���D��a��<�Ӽ&|�3� �P��)��� N��'�MԌc$�g/iڒ��Gg�M�6��tvN�ԃ8�����A�8d�s�yTTU���b[+j
�'6�o�W�ӝ�����'�RnZ2.6M���$uyq鞯��0_������rK��߹���i��'�	� K��Y�H�Jdo���q�q�*��74����2���]5䭰�s'�8Uz\N��\�`NЏ?��1�I.Ն���3�`��%s����)����ݝ�Z�������nԖ]��q	���RN^��;Ym����o��#�6L��	0>ƀ���)��D�{�!0��@�]��)LM���
�I�)M9��d������ڂ���<��PD_��ҹ��7��Ci�eI��j�2{�� LI������\��`�h�ڞ�/��S�t�8ulp��q����@�O�wW��R��<�A����u����ӼI.�����&� ����� ������;;�����y���$�;Z�wQ*]\^S/Dܘ�ԍFd[*H�62s����`"��)~2%��#\`�*���V.��%F>�. �A���=�Oc� נ���T�g֣������6��6�WP�/�FU�X,!�����AQq.;A5J�ؗ�~��z:`�*_/ה��DKi�mt����܉�y#[F����t��l�<��)��N��~6��JӨ{;�a͔��u��r����e!��ӳ�t%pt-��a[�Ǽ��~"Q�<���ppQc������/|(�>ֱC)�����hh��d���]\���oܖ��x�OMz̉��S&���i��x>�G�֊����@Rn3�f0��}<�K�}�'������h�laK�����ݫN�L�R�$�FF�K38�9�؄��@�Uʽ/�V��A�N�)�����o]��_�\���4�UI����e�t��A;[fIxSz/aІZ��`�1��o����ǿ+�;KՐ�ع}r�ٰW�����}�������c�e&D��Sw{42����� �!!ۊ�t�����=q��X�U�
 �3��ʕ��~u���$�V��i��m�nQ�����27K���έ�~5�m���zp�5u�78�� �.��J�&Y�N�X$�hluʳ�-1�]$�����W��酋SuԸl�n���:E���R��(n��_j���SS�c�kƧ��=�9S�W��!�u��V�7H�% hҟ<0�t�˙�������)/y ��aם��t+�
�5=�k��|­[ c�`�g�[~�p��f�2���K�Lh�������Q�&94
C��r,���Hμ����"	f/���'s8N���,�dd���>l��̄�G*����_�xK)��������({��E �31�~�Aː�#9.(�?)�
*̻q�=u�6K�I5���)i4��l�ˀR�\C�Q.��}��J��j�k�|
�oW{r�vcp��0��s�U|}�}og�������A#�(iڌ��ދ�2_�Ђ/r33H��$�ߓ�
�z�*�wiDb�f=f�*�ϰ���X��~�BU�<��[�K�P\s)n��O���:GH�v��q�(�/�����ur�v-�Ǣ%��g�d+x;�Nr3"�7��ut�*MU��m|4}4[B	����2�E�>]�	4�-v�J�1V�w
с{��D���	�$p�qxC�'n�v�%8}��|T��ܺ(�v�;9b�N�#�2�.J������
�Z��x��>ߒ�x��L����~��J������dZ�p ���<�h3����۞`O�����r?�_Xx���n��Ǥ+�*������!6�a_G���ͳ�{�Y�;�3������s���w����!`S[
���o%ګ�t�(�F�O���4�G-9|\cIk,�d���rum�E'I�Ც���V�҆�D���2ĿN6�2���V�;�1u��b {W���(�~�3�ǵ�A/RKY%w/|Iٍ1/\�zly�[�h����/i��Q'��tͼ�GUu�tz�.��B%Q�g��xf�������0M��v�G
���p�Cs��1���t��9{����.��1��D	�e�_)�>�q���_~"��2S@�̈�׾�n׹]h�2	��V�3ҽ���/S4�'. k.3�L�RXV�B��*
�m<��D>h)��3�_�刭
е�|ǴP�z�·�w���9D2�W1b�vZ����ۼ��&�?�--������*Cz]��ZBmF2y����X�X^0.<�`���-�c?��˹�P�W�j���-�3�P���J���.��,���K@.=��Hx$�1VZD#AOC��0ϫ3�,�gy:(_����I�[��y��,Bۢ�azr�uY���5g���2>���+�|K ��O� �[$��.��{�v�Av:]�,0J�e���+�bSEK���4-���e�@�/Q��1�m=Hb�UAmz/X��u�Z=<G�1 ����, ~�Ѝ��ߏ%8ߢ�v��Y�Ue��
5�A�b�g��ҹ�0���Vّ�6�"<�/�;����:����͝��S:�L�2����*s:�>La4����v$����z+<.e0�ńk�yg7kw�6O{Q�3,�u�h���H��n�M�gs���#�=C
i?���`?5?!^���}ξ����7���,�J�=q|dz�Qf2m��`��A;ֈB
�Gp�Űn��|sA/|��QQ��^ҳ�Zzȑ���,R���|\~��)5���4��%�Z��5��\|�^"b�}H>?���Y�\b4R�!�K'�����W$Ho�kj5:�����9�7�h\�8$6S�z\���*���[��XۚƮ��!�w�%y���η��q�`�y�u���M�B�~`Y���Ou�~If2P�sUo�sAܶ�B��%#��+�vvQ��H�Lˏ1o��� ���E�״�����V���x����y�%��P���b����3����թ�����m����g�6���24�L�r�G��u��*���˸�Im�b|��C�v�E6���c�D�6�3�S%�����̦ͫ�ʏ��K�~ɩ��E�S�j�W{Gk���u�BC�;5Y|��z�I�T?��5�+�-��J�C�$}��=Z1�髞-kN���BqW��-<��*`)H�%(�_3+'��X�p���`�J�0��h�jW ��l�H[Uj��=�� u8���b���!}Oǚ�3d�	~�!.M.��?�#D#�O]}�6S�ֱG�Rm,�3ac��	WY��rܘi��T8N�>�ˇKy����o���/<�zz��~>�
F����@�#`b������X�)5ݐ��Xn�n�eb%LYť�3��eGV�6Yt]e�}�u{� '�>�ߨ�:-����9;�6O�{�o��3ژ�m���Q�Q~����*��:^���mx�;���#o�Tc����
�����>b�}8FoN�s7��>H(d�Q���8#0���t���V���t�rBm��K�t�� �F\��w��-�G%��	�e��[�Ƃ�jP.@�5���k^��3�(�����ٹc���{�VϹ�"�23�p��e�0l1��W6_��x/p�C�����]�@=18��{{G�'"b%ׁ��-�fa�5vЋ_��1/���P�z
"hQU_�4Za,��'^�Y�״]�ca�PL7�,q��z�}z�c�@`:n�9>�3y����&?��ϲ�����9�Q%h��I�z��0��h �o��*|9�/��}��8�5��,^�Z�d�f�(�Dk�wm�9�$(���5��]���EV��S�;��@����v��Eo�B���5�';a�-�K���׷%.��w�G�d���$H�2j)�;w��߫#M��\>�j4�۽�d|����\�P���&�업ؚ��
�2n��p~�_��������|5H�s��i=b/�B�+�}/x�9"f��k�cO8D�))���/1�������v!{R�Ju��	T�*~�.�N�^8�E\���VqS}[�WH���ѡ��W�\��T�����$����ӉKdJ���w����1���J">c~�����"P]b�'�/�V�����$z c�]8S�\I�s����>u�N"����
7�vn�ថ:ő��nW� �i�_B
xt���E��}�F��/&G�i��^�&Q��`j% �&��4�W��aX�ݻj�޷�oY����`����
�l�s��#��f_;�w.��.�aeW�O�	��Hel����Q?7�j��E�����!>�G ���\TC�Tն~������V�����"ga���d����� �w�+'�4�p����.��wƇ��"Vs~v>:��o0r�EMf"�C���F:��$��z�J�)*���-,t���N'!���S;���5�!�/��c����XC�w�Ř���hkRի�Iz��/�:DD��f�/��ll/����b�X4�v�LL�m�E�9�_���M�����Q@�31[��s�r���ЪVl�����Rp9�!IT�q��wX��Q�nez}ě$e=)s�k���uX�}9#K��i��K��d�=���j+l�SGe�v��f���P�b�q|��cR��_��8�.�E�G�$�5r��U�j�?���ϋ�S�����J���6wϮ���.Y/O�a�c@��I-�Y��w6翑�k&��`�=�gf;τW�5d��k���Ǜpw��œ/���_ͅ�<�|uH�;���_���ಷ�/WX)�U���ۉ����Q��l�-I
2�1���ѯG���d2��F����	S �tٰ�����єJ��hE�)�f�������z`X�T[)�"�%n8�_}L�Cze9ݠ��`$��H���}�z�d¯��������������JЖ�e��ʒ./y��V��Ms&0�
�;z���QÃ��ԯq=x,�@˳C�/�l���1�W/ck ��n�)^�v[�~��h@@j�v�����!R�P��|�W37qKq]���B>�w�l="[�]��E�3��Se���M��ncái�\����k����V��<`z-E��T��D�_(`����R%(�(��K6�.�H�	`��8�
KV��"/����W�����ɾ�!t�`��&��0�-\�Xǒҕ���dLBg��m��
n$�c�2B�U0c[�+�d5]�`����w$ݗV�sH�1A�me��Θl�&OG~΀0�8:y̫7L�"d!)�pY��E�Iu�&\����ɰ1e�Ө¿�'�ĺ��A��&w�t���h��O~����1)Ő���K�������h��Ѽ��t�B�S".sB]����X_&����J���8RLF'�[/��=��,2��@�tPH�ż��ܓ�D��e�aZu|V��L�|�t�}��w"t�}���ObB�籑��[��z��o,v���a#���^J�MDtet�>>ߺp$⨌q�Yx������7{B�!xAk���Rк&���pZ���|ɮ��{L�bď�=f�����
���xNwUjz�F�hP7�gQn[��gC����㨫o��/D0L���Pd|����?��m�r���Ye����@��㫵/�v���%Ѻ)��4�s�w��8�Ըɸ�
��q��.�����x]���:S�;{�F&�U�  v�a������Ay���X�t�q�YAM�ۅȕyr�����豾�� m� ���:�^�H�V��H[���"����s�K�d���墭/�?A������7<J]��6��r��yh*�~xs-r��F�0�l=��5�M��[�Ji�ogx	�c��ȹ��2�4[_l�Q�>�ei�(u�C�$��?|��Z��X�Y<��B'Xg#�M�^wrF�Qžx���.�.&����?>�~�`�b�"��P{,{i� ��b�ܼt�ұ��G�N��t�`�g���7�7|T�"��_�U�}z�_6�����x/;�;mȘ�X��y�n�Te($VI��y�G�m;|A��[� ��^7UlKA���=F�Bu�*�TYLam`���Έ���3k����XUC�mY	�����gb��t���8qsi��[���ɖ#!dMl�W���Im�i��m�Nߓ/$LC���	s�U]+��yGvM2d ���nۺos�?�W�s����?�A��8�ޭ9�����.^�b߭˒_��	`���Uǎ�uZ���w��N{��2�S;s��F�Y�Z���אg|	������J9��ϝD-9䔔I7+U�r�]����="�c�q�w�&�b��	$iֆ�u�Z�*ǻ���\:��Z{���S�.��x�.�j�GBl��M:���whb�+kqx�Mn�fs�x͐�p	��q�@%�\��*�፞{4�\���t{�,����@Tk�?Fǈ.������ .���0� ��� ��I5$z�Iš$���uu�8�I�FG��-�@��mY��;���������N7*�r�1�N*{�Xn�"N���5'U�⏖��a6�����2�<���Q�&|.��I��P�D�� �ݖ�+�f(����7�X��
�p��R�U~S�F�PR���\�KDV�0�ܰ�����r[#�ۈn-�����/�\����D�
/ni�>e` �|�Y!ieZ%��`�,�b�K���?]N��{�\����:��C��c�{X.��>�m����#�w��l��ܗP4�H�2&�8c�j����n"�ퟌ��#����ݘ��G<a�{S騐Ӱe+��V�z��/�}t��_��8މ��p�
ry�z�}������m�n���ט��^���HO�/7�����ߞ9zTtj��x����̛Cz���}�}w=v��
)K���%
��V�7�ĮL�e��}�4���h;ҙ�n�<��Ɠg?��p6���{H�h��N^^
�N��G7�I\�?l�vF&�e��pUuO�)�i_�Ɍ�7_��/Q�� �~��{�z�t��>�YoE�wD/���QЫ���:o$
��U�-ԕ����W�{��l!M���e/
��������综�ܿ�-�V��(x���u�af0o�ioj���Acr�_n3X=��;4�x}�rTH���m0|�>q��{Q3��]�`6�@�������t�B�V{%AT�A�r��6�`�ASGE��A�G������j��Go�!���`�2�n�|�%�d���_���K����(�y°�Ի�Cy��R'�����E)e��� OB�=)���k�MO�b.������7�� )�Cҭa�`D��&U��vo�{j�;��ހߣ��Q�����z5�3+�/������7F;�W�Pg�q.IU��9V���Dgq3�����B�֭�o��g��;�+�̈́����@���B7�������{:|O��)
-�~�!:��5^��O�������(Aŷ���S���W�(�/��p,��J�T 5L;��D����P]�kGҤ|�5�ߞoyP�'Q�=K-�9�N�,�I�}�Dy!~KxEj��x�#��gIDӑമ�*P����%�P<3���+��P��e���f�kl��ߵ8�U/ԓ}(�8��\���:!�|�H�A�ԖV��E:�DG���ڑ3Y�׆�K�
Uf!=��=�Fƹ:����
Z\�=X��;O�����6�.��E�+��UF����� �({�����\1o]�d�����i��F�BO#絛m�}����5�.�h�Ŝ��4=���O۞RG�`L�I��Sh��Pǭ<�yF�ј[��ˏ�����$���	w�5m�*�}~��Sj�5
fN~��O{A���Ր �g����o`u�%#?I�) ���
��U�2���У[�����8n̮H��M����m�^'U�(O][�'۲�+(�lb�l=&��
�l(
��e��{t�F�&�G��q���I���N�ٖ��j��c�@��-�ZJ��d���'\X��T00��}~��׮)���1�V��s|�q�E]r�	=(�7Yc�X�%����X�~49}�d�{!�et76(���	nخ���]yC���5�Ջe?_ �%n��Fe�����Eʿ�O�G��l�V��.od�M�x���4:f�GN���A�wꟸ�rS/��Ew�tK���}����n�k��OrT��?�tF���%����1�tod)�����:TC� =���d����8-:��=�?\����>?�;*����jN��kĩؠ��1�|0�j����wwX�>>` dV\��-���HE/&�"v��mt��q;ݤ<̄�?�$�з��?�+��0J��w~DGaP-��R�]Ӛ����Z���H�_%��v�vZ!E��֮��S��]b�]�'�V����Q�����"���Tb��Qi/Oѭ1�&s��~១� ��a9��s�2=�rVU�z��؄�������O'R7��.ؔx�u�����䤝��;H�iX{�w��"�k��r����T����!�0Q�k[	D��#��Ѩ.TV�8�������˘w�#)Ss�d�o��}��4��ޅ��&�<49T��y��Ӧ:u_�P2�����c��b�Ԛ>�]u�H�OR��JQ�5��3�ȻoE�qHF���ez��F*㌆n�^q�$��V������!��:C�;aN8NX��Ɨ&=4x�-Y���z��k�\�Q��ڻ��ߞ
h��W14"��J̱���r��L_�����@���L���f���jJ����g����>��ؿT�}�ə8�/�<�6Y�,��*�;�9s���{$���6	���

X{8/%��f߬9��:����t]��i�zwj�T|:�I�1~{w�ف+�8�h2�������5C�2^MʠtN����5�8UP�m��Z�Z��2zQ��G|�cݧ٧7�وQeƍ3�No�B����*��S�2�V��NYh%Xyv<�A��GKq�sm�;;qAےb�;�H���Kd�����O�W/*/^�,|�;�<�cT�u���������%�3�3\W�w�m�U�Q�x6	M���Z��
Ը���t]��M�t�k��E�1p*�3�;5� �|��Zl�����X�����'���=�N�,����>f�)�� [K�� W�Q��s�:[�(�b~ʛ�ߩCH#�6jO�׺�X�JH�$wLiBAi�����/b9a���=.
D1{|�ۓ���ǵ�2�P*���=��J���_`�����c��0G2�$766F4*�2����?���v��G������4���ci�m��(ME�g�苇�ΆP�DA����!�4�h4���6Dx;}�U�I�����1��S��fn�e�U��}�K��тKk�R���ҝ��P#Nq�וgʮg�� 9���ʊz3C9P�@��ӎ��������I��o�a���|F�p#�2.�m�O�K
���k)�{�^�H�#Gq��Ϲ}�>�L�/�����Ƣx�Õ.E4�|VN,�PeS�!�~�L���u�r���l��B��5�_'Q���+��6�e�� �[1��D����i�T|�1@*��|j�S@�Pv�a��QE@� ��:rq�B����*g�tzhZ�>�d�\&y	��0�8(�w���Z��<t�5�,T�d��%f ���|�M�
�D�$� Ŗ����BCC���Z�	��B���.��*R�2�P���/+�����^�o�#g�Tl
X۩���{Z�I	 �vPN)���^Iӽ�Y��C�f�c��1e��z�" HK��@ā����k��c� B�N�����l��I8�N׬�a�LGV�JE��q̀�F��̏�u��O�1�C۽O�qW��sWP��S�'�q~��ڲ����[�H�o�Ķ��2���~�p�JV��g�|��m��.�9��m���*v�e���|�&���O$�v`>0��æ��h�c���$D�?�&b�D��fV�]Ne�5\���yS���vC���)N]4���v|�����+osQ/�l��$�{���tI�y��O�W�Rʀ4�r�R��RR�FSѾF���'���sv#��'�����faqȄ�#N%D6:�cz�Y[�����)��	�E
a�!�7�J>r~\�b�G�n0i$V��yk�W��*{���E6�"��z��_ya9�?����T8��>�ןf�~8���x=�g9��Y��0[\F'4�TZ�@�ϮV�������,ӆ���B9Z�iuf��~+�v	�
2d�md�T��zA�Խ�6���W:"����S�,%�:����j͆A����w�T%z�Sc--�z���|נ�a�ӵ�Kj���Rbk������G	�����s2_���>U���~�f��l+:��v�(�S��Ҵ�����!v��\T&���������&��B��- �犂"	Ty1�c7��o��<U�r�ṡ�����s�"kՍ҂u��T~mW�]!xу��c�u����}���*��=�&#q��/kVT,펗�Zݡۗ���N�K_eĝe�,ɲ��w�;�381��-d���;�~��A^߳v�䬛�έ���Ͽ�Qսp���nL���/f(���2����%P��SE�߲)S��ӗ5�5r�m����^���ۼ�o�[�q�x� }���y��f�%�b�e~�X۠zգz����C*�,]�!Rq4�Ot��?��8��wC<1�Ҟ��vߋ�����$Jp���J��Kd�̛)�o(�k�����YRe:�1�< +q��U/�[pd��ɶ��~�O�k��F+����/p+u�������)�� 6��~���g��g��O[�xĩ*��d�@3�Z�O[�T%v2
�2e�W^P�mv����AE'Q��9�%��c�U
8º��u����Tj
��^s�}���0�F����,��yk�9�������i��|~��)�b9i.��i~mYX<�@ʽ'�g�ڰ��,/��t��uH4�t�6�dMnlKy��LRb�5���[�h�>�8�S`��T�QJ~�&������A�M]�Y��wI����GL��>�*��h�^���1MWg����h�	��n��3�o$|�����w教���U^j@[7ӆ8QB*<R�I�h����ns�S~ym	�7�K��4$(�|D��[����=;:�u����~�7x��*��sޕ����B��y�3V�KTX�˗���N#^U*d6"'&�my�0���3�E|�/���a�Gﭭ\l0`�͒�����Z�&E�xeKX�z���;�X,(����r���<E�i�Ӂ�\�����_�2g(6
m��E,�������iUa��U+��x�X-��	LD%�!e��AG�	C�A��X��4�Cɓ���/7�X"6�����t�/��^#��\�9���M�6�>5�9"BT^�(*�i����8^���Ԣ�����>��wB��r��*�zϗh�S��~6�K�OV����K�Qd��ԭG��O���G�o`^�=#+Mz��E#�x�!��<���w��(vc>�>��P#��!A�[�΋�5�薯�\ .��_��9\�Zia�f?����Xr�ü0����(�p*״D�'�Qw����7�dW�W�T!�ep�Ѻ�5-��Te�
ڵ:�Q�ן	�������;��d%
����ˎmb�<��Մ�� �a��#|gw_�ޟ<l<�Do������zw[�M��=�{5�=rԉm|rYzɳ�-�{�+�o�C�\2�b��y�/�!��^H�5a�C���8����5dP7Ԥ�F����4;T��U 3U 9�����60�=�_��?/[�`�tMو�Ǭ]�S�������f}!�It�.ъ���.�����S��Tt�\�O��k���t�3&`����D.��0y"c^�K꜑���`sK��վ��W�]�_j�v�mԶ�g*{g�(F����[V{��尢k@�9�7S��N��>l�=^A���њ����#�PD�	O�T
�(��v!+�'�g����$���IC�[(c(c�;?$~$ڥ �p���rKT�1(�5�)>gU#��ӦAY��銡�:�4i�K����J�Ê��:7B�F�	�1^����{�ܨ_�&��x"��"��֔߽7e���N��C� �M�S+��pk�xG���rE4����ha/7�C]���ea��Ca%��d'R�F5-����CqjO�Љ�t~����iztr��,ƄiW��(mC6�m�I�w�	�%��;��X�x�q�3�e"�5P���H�ӯ�����q̼ܫ��Q�o�J��[~���q��d~�E��~�]zNLN�D��%��F�PA�h�
"�[�l�,J�N�<JNk �!g����1.s/�P��$��VBwJ��v�,.�0��?�_N��rr�]��ml�i,/�9b��B7�1�,=I��vY��Di��_J�C�q�x���������_�dd����W�K5�A�t[4�����ى�n�>vƎiJ[5a���*��s�0;�7�ae�����E����Ǻf[�_�C����������aƏ�5T7�B�B���l]b����.֯� .*�)�I���Cl��>�;52o�X�SN-ټ��@%:�U�J��,d�_5�*�_���S���*t=(:ȸđ9P�c�.+%�ME)��Q^H�պ�wl���+^��c�!A,`Ў�"`7n߳g1��z�!��hJҮ<Y枿�{�#"/�v{*�w�\��JN����$�{d)7jd�o�hf������*�4&�/���`����%�oo�w\-+�]�@�zu��-	�c�//v�,	�������n��ʬs��ӡ��NCo�=-�XQfNz�����,�n_���Jev ��a�x��)����D��0
�cl��j�ۯ��G�~�c]��m]��I\1n)��k�?�Q��Ĝ��ٺ��P�VIm_�j�N2:�+��0U�gR�;�(?�a�ރR2u���,�Rgp�POZK�Ȱu��M�^6]%���l�g�K��q0A{��/[-���45fl�x����>}By_��!��ݸ�{�C֠GF�!����I2�6;��J����$��,'g^ʍ�HGU�@�Y�!���R3�a��8�]�9���C�
�v��|7��w�hxd�_���x����y�x�`��R�˩������Y��gvW��M�"ل�N'���ڨz���&���LS��|��Cd�
}��pՁ���qD�d��銘������""�xs��Ӣ"��_����E��Jx�{
Gs�[�\��5�� r)?���ZlV=��u�=����*rI�b-؋���3[�{��<x�[L�1v�_O�����l���\EU1}����� ���^Y���}xXx��U�9c�41�;�Xm�h��\����L.�&x��v�-�)l�e��m��2RE*�(v�XP�8~�4��ɘ��Q1��3�6+A�%�N4����GJ��ws�Y�j������1��+��Ҡ;{߹/���<�Wf����S��^��4t��U�c�G|��+բQ'gV9��V�ʢ>�csû�>v��T�P����>�����w�P���Հ�`P��+o�c-*�:6D����?~�Ċ�.��W�S��遂�0�i��%#e���"Z��]�(�I;���"�fF�]5��]�7\o�P��sr��N[2��#l,Yh�"�5�%�@l b�d����O�^���6M�6�m�hr�4�m�Ic�Ķ�XN��<�m�i��o�y�ߜ��53kݟ=�Z���4��ad��~��͆7�tU���r�~$�Adx�aS�pb"�-����������#k
㇍��b��*�q�*�n�a����:@�d�Z(2~䰅^�$i���^�S�%�J�,�2߁ds�������5FW�?fO�ʕ:!�ΰ�}4T�t�G9�>l
WP)+��~�Ň�ɫ  HP�*�r���?�D���M��A��!�4뫲�m,DHN3���#��C�+�;	`E����P�N�U3М�~�������Y���[����M:�֣v���>�	���hT��q�b�ܼex/3D��6�;$M���-��tim�_:�O���=÷�8�;��x��ޏ+U�W|�3�����C�`��B���r�Qm���Meނ�S���E�\�$Kj�EaUL�]p$��)���P�Eej2C)#�U4F�.봠�=F��FScSHA!��s����������H�nЭyL,���a��G"e�I�XFc��2�����|�1���%g�9G�A
-8��R�ܢ7��V� 1��u�p[��e��׭=m�n|Z��0�U2�M/�uE��exv�:; S�`e��h���U�9�_� �)A�^6c�X�����K���G2�0Fc��r⇹�tk�6��N��8��1��*x�O7�����ϑ�>����x\n}NF�0����?T�g *�����9b���&��`����"���q]�L>�����!�}� 38.H��a���ωc}����fe�#	{���6,���U�l���n3�f6��u7*&r���,>NG�Q�U(v�5�E��Y4�{���y<��N^�PW��.:3�sc}3a�v�	�k�^�!�MH-kL���������S����)VD��������������r��V0XX��k}L����*�Ŀ]@8��k:nW���C-�Պxt��GkX����h������Ĥ��cNK�6�3/�%���f��T����-�N��xGS<� �`�(�-}�;���^�Y�aΰ�����?�r`-�Rt�Ͼ��d�kk���$���1s����	���5�W┑Ӭh��r@�Bi%r�è\��yz���>�E1����Y�h����f�+�-�-a!_�����	�%L�|L������c"�A��)����Y������a�dN�>Q�qA�teyV9
��\�{F�quYY�����[��� �Y>�_��r���Q�V��
�!�=�-���LC;��֫�P����O����X�pL�C~�˾���w��$j9$�U�q���N�7t;�l�,�y��t-c��s-b.e��� ׬�ĭ��ڀ���ẓv��r�}�[xס���������^���wϸ�k�-eG�!3�Zv�����Ŝ|������6�?��V7�ގ6i���.����Yga��9�ѿ���s��
Mi^��h���|�3���K���-F����ڍ�����N)���4+T�(y�5��&�0wSVnc1�C�HQ��/���þ �f�c'.���Ŵq׽bCc���b192$��H�CXB��I�HP��4?+^X� kz��������m�\A�#�K�b����V��9E��ʔ����<c�wN�ί�E��[R2U���S֦;ö�L�Ǔ�$�o:��T��I��'ʏ:�=1��p����Th�c�q�?07>SyC��2�	|�s\!~���3���V��V^��uR��.O��r�kU5Mz���'�lOK/O�x�۱�B��Q��0�A�{�<\���o�I�ӂ��]���N���9*4+�s�8b�c�ܵٴ�_�[ �T������Vl4ɮd��j�������k_�ӧ�����usl�k�q�Fe1
�-�1��Y2zL�R���G2��w�;����^{�"���������N?4R��D�H�&���N%�c�Q�y��:��gm�B۷yk2αW�	d�5�|ܮ��;S�x�z���I�DU���h��'��n\{w��3��9*�������k����G�	k��5�����s��Ġ��m��m����M�ΐ.��"ҫq �:"z��Ǐ�w~s�XŹ�B�Z�L9㋺���>*�Z�93�u>�WCq"ft7L�5�x��U�� ���U���_�#cڮ���q��r��!��*Ku"�Jv;Ҫ�F�<�']yq���(��#�ҿE\���>���� �~i�])l�.N$�����l�~�px|+D�m;QN��S�o����ޜ�0��dݢ]��}j�T��n_S{�����bC����w�6�Fu���[t�_�1��e��9���`��
I���ҙ�O��l��ZԺ#�JR�;�Q:J��X�T�.T#�&c��� �~������6�׫���}=�m�E�Yg���T��t��nL�:�����?��D]qR�8�tЋ�N&-��7%�G���q��ّEP�;v�e���Ӵy�� _uZ !vg,�د1s���1�f�y��Jy�U?�.���yQ�	u���^yq�����}�&>�t갍�,A����|����Z����H]��i/(���|����|����0�owж5���Mx*2�C�l=��Z	�t�J�o�<e�X��bӠ�
�D�4�|�x��]"_�Z\�^76�t���6�Ő�,ڮSF��jt������V�����x�ӓ��Ec���+z���[S�`�������p��Ӯn��a��qɶ��!�j�'�ZϤ!��}��|����~��7O�V��6�r\	�R�d���w�Y�C���|�
1�Y>�l�W[���ˬ����ݪa����D�L�@uN��`� �c��Q�2	3뗾�$k
3��ʆ}�� ]��t�NNB~�~�/�f�U�
���n��I�*̗�Z���$vѦP��ڡ�x�*��=��A���{r�F��s�����\���%2�{+�IYyz��=�.F�<�鞼��&��D�š+���Y�G|Ցw����>[��9D�x
Q��h�1���4�0k6���w?���d�r�6�Jv�BƎ	ș<Z��#��|=f��@��r{��}��7;%��}��N��,'��{]�+O�/
	���Ϛ*io��T�=$�{�~]�v��\��k�\�p4���/m�������n���(i�?P�*�L����0W?��N�7�o6]�>��o~�^�~p���/'�N��\ܛ���u���_N"B�$t$��P�֔��~���#D��B��Ba{�)G�CH�[	e�
>������ c���ُ����C�E��� e�K�D*:C�5��uea��'o����<�u0M�D�@�xkp�M�%9w�r�7F��IKi�en���,�\���F�u�w�d��"V~T��H�hwW���_wp]/xt0�K��^N���0���X�bz߯����szNu�|��ak	s�r�����y(�x���AV?���Ag��T@�]}T)�U.PY��'��"�u���M��*`rM�]zg�Ԑm4�m#�K����`M�5:��v���� ҁ5n���Q���0\����
j�e=���D�2x�K�d3��xL�����-2����xRg�}�Ӂ-�gF<��û ��8���#��ß9�/jQ{>\�Q�$Ҿ�����l��7��-�m���ં�}~*x��1�@����J}8(��
LxƪIh�ƞV.M;z`ֵ:1�#�
5�^XA9ML�R�(��[�a�IT�������`�I���;f��B��ے�Xߦ�Y������y���"-�v���~��P�N����µ� 1���b�j�o~$8�)uz���~���C�t�׌&��WXHP�D��D�6�d�w#��� �<Az�,�հ��|�����`zqPD�;ؽ��ᆸ�>7�47yv�IӋ���f�-���Ȇ��2���X=�Qd~�/)q�5��Q1�� v�`��|��
c���O�W�A�26�ԧ��~�Y�I�{%�m�&+Z��w8�������~�)�_����DO!3e\G��pJ��<4�F\Z�F�I�0C)�X�5�h��5j<Io|�1��hߥ��d�A򈷙ɮ �E�E>�X?Ke�Kb����0\�0yK��'�%���{5�F��%�-,z���x�3e�¢�m��S�`�I��aݩ�wa#{y$�Gx�&wyO�/_xk��[�s1��na�8"��%�>d.8��	<G�����V���!��t�d}����^�c/b9yDOF@*��N���^��@�"�Q�g`�d�@��9�гV�����]��l'v����r�#�I�>�����R\T�+k���Bޱ�O�e���a����S	��9T�A!H�c��䠡��Ŵ��C"��#*$�@<�ּ�n�V����A�K|}p�&NϝOUq�쌜�N���#W�S\Km��9k�E 3$[��Ց}TD�I֏��*��M��,��Z�q�"���S�@���ߟ��A�u�l��mh���Q;2r9�2,��Op�������j�e��B�V)��9���H�;���ŀ�0�K��a2+F�9Ɇ�+G���pҧ����<s�^gu�Y�h�Hue%�"���<ޯ}#t��,Hm��eݟ�z2�g͖��4���Q���?�r(�3��w�㜚�C�k^ß�K�W~y������>7,��pvٺ�c�4��6�`x��RTqr�uP9�c]��y��l?(�Os"���`�����[�8�XVZ�;����ldOn;��!��HfVk�܉��}�׶n�B$�v����k��*_�x��<��k����n��`1!8IK�O$ɗ'Oa1�����3=���@����Akju�AV:f9$,��'�J��3���@��N*Aw�F\�tsc!�j�	��u�/;�C��7�6*�Ҥ�+0h� W�p����D����=?#�4�ٻ6" q�`j� �h�	�bF"ɐV��#�8��H]A��OB���WJ�a��2v_R�#n| tޚ�65bɦiZ{fl�̹�_�̮��,�>g���!�����D��y6Q1�	W!�.f�0����r��F����� 9N�<�����#�y��ѣ�<��1S��� X�u�Ү�x��$2���t~��l�I�E�C��!G�?6��$��Ր�a՚��M�Ⱦd��J����m�	�d�hҰT��Ls�җ�/�eVD��ma<ur���� pי�L�,?���'7-].6�P���I@[�G�����0T���1��w�9���q	����ֵ��gAf�U6�g�--'�h�ܫO�5��	�
xR8d���)Vt�鿱�J!�����£��~�r�}�ƲB�!�������4�p�A1@?�^���V=3������ŨЭ�l�K+�D�J"�������AݍQ<�DRr�S�'�|�IR @b�s<��DA�M�v.�9QA�m������aR]ty��bB|�q �Ԣ�����/��	�<*�8���y8��S��Q��Wp"��Lᖏ4�����Vq!!V��B�q,1�*����g��(����j� �ro%)v%g����8g,���]09D��s���n~D�댰��7��o�t{��Z�d����"�ꌪ�V3��^m���r�n`?�t$a����;�A�@��{]��"{��(���6�".	%5d:\�Z^LLNL�$R��E9��mu��� ��Z��]�-Mon��L�H��=���BbUD�2�i��yA��#f�"�y�&<�c7����8�O; ��>A���צ���	���r�����9X�K+|[�^�ˇ��=�_��/�6����w��ݛ.��q~�on\;#{M����?�_y\fh�������<]�ty�@�$s����)}x�/�%�s�>�_h����.���>5?2>O��z׼>	<���J'��]�"<��9��<���<���Y��V�)��Yr���^�l�광�t�Ʉa���S���?GNG�:U	��9f=	D/�(����SL�Bg�����a^𬋄ǧ�;s@��ϥ�1a�A}��״�́IñF#D�L��ȯm&�߿q����t�]����#��6��z�N�`1lAqɂ� "u�	]$��۬�V�b_��o��s�ה?���38�P����;��(��m�b��f�����p �$}��H-��td��D�Љ.��?������3u�r��<?5e���03 D�e�3m�\o���S�7��p`�~�B�͈�t�y�kj�i���(�4q83�$rf��'R�ehW�z����f٪8�oK��Q8\���!N�>8>�_|����Δ���g�+�5a"�T�%S�7>j�g�ah�Rхh����//�i`���C��!2yJ���x��3{��Z�[&Z���#����@�R��+���s���pG����t�uZ�}\Ւ�ˮ�gS���'0I'>�b�&�<�z�ycef�:�MV�]C���ɓ��+�3���PҁB�b�9��GX��i�mQk,�Ø��-0W�𣏕�˶"�Q��4eꈚ�󖅂���>�<���
C��b&��g�9z�kK7Z���cq�!�!���f��.�GT٤$a!���ߢ@�=w,	�ᣣs�[�����5��L���HΕ��p�9��|�JM�_�/�J�\���\�)%�<����`���粶<�b�; ������R�]l�z�z��d,)�y�0�E����щc�+[�����X**�8
4L�5�"y�����F�\��fi���n�zv����)R�#h�"ˢ.��䨉��e�A���N�&+�_F�dd�BƭdJ�*N�*s��)�W�;����2��>�b/���}��ǆu�-t�e�F{�G������YL*�̡_wD`t��	<�]���G��LS  �\1e%�$4�m����.�;Tr~�z�L�^6{-o��+�/�~=��F�>5ޮ{�7����0��9ŷ���n����Q�,K��f���U$�rrָ��%��[k��/�}x
���D��ۗm;��{��M��p�D�3Z�r0��H{KO��.�H#�vH�~�PF"%�΁/5�ǘ���)���9n|�9ջ�H�YI������[��#kkT�p'-������@�%���辐�$1vk3/ gD	�����N���7�(W_�CA.h�Ң��]��jm�^�5l;TLmT��'*���є��6�ĩ=��_�I���<^ۻFLS+sw�ZE��E��Cv��8&!m�Pe}Un�sB%J�	ZNw�[b��(�H�Fk77S�WW��=�����򲔎ݵǤcF^4�Ec��/��j�l[;���M#>�@�@W�N��Z��Ǖq��J5�q��~ q�S����w��j�~j�����p�@��
���_fU+jY�ܚ;��´����RQ`o�RP�ڱ�6��n^��&�&�_@X���;9
^��JWy�u�]X랲ݤŗ�0�q���{�2�5�Ŭ�I4�&���J���` _V��I�,�JW����M�-)U|E��,c����'OR�d|�lU�R�v.��GF���p�1';+�e~�o�0A��+�s�>���W��8�X�GvqB¢b.i�*�{�sp3c�Z��S��r˦�M$+�F؉/v�P1�ތ���0�x�����P������k�[l�g9Pp��	��!'=0�q!339�`G���"D~�����xUعT*@P�D�*�j���.�*l�N�	�j�O��j
��V�쁒k)K�Leն��1��V�b�d�U뷣�H��h�u���"[�N�I�+H��d湔�q������6�
��g�6N40=?o/�l�ót6�`�0�܊�/��������.��E�}��K_u��v���)G�N�'y\4G��_Q�OA�XJqɔ��E��XRc�Q���o?��̜"���w������ �� ��Mn�{�buM���������{3�ޑF���v��L��S�IS����3n�u��=S��uPF�~T\�j�{�>�tC�f�E�1���`d�CLӺNK��0-��kr�dq�K�iu���"޼�X>��JFu|5��kYp�N�����ɮ��[/^���Ո��#�`��Xƴ}�]�����@1i��r��t��`��G��%�y<�U >þ1���.�VDAe8�g8����fo" ��hc~��?�1y���By�31�?g �⯧h/�$4^�+�����Wj"d��8������Yp��U���������:��(씃*�=��R��լ��8m~`_�I�RBf��0-�L�1���/�<�u����J��f�����bEr�@�q;|�ٷc��lnO��3�Z݋������12��Sa��A��!�GǞ����ك�2L$�NJ^�Ķ�5���x}գ��C0�QATA�Fʆp�.��.Y�JL�_�LT	�)#[%��oX��Ý	����}���ӹ]x�1���H����y YtM�φ��L9ɖ�
���b��z���$�"�G+^Jp@)�B	S��We�R�����"�R��ڜ'ubU���,=t���:O�r �'pe�p{���д@��o؅���p��F�E�k\��L���_� +�:����v]�m�'����M
�6��+����g�r���(M�`nBٍTt]�+��*�$--�;�KoG����4�&'2��Ox�t�7��������T����k,�ö���o�U�l|}{�1�;GqL1�(��$V�϶!���X{��>k>�K��펵v��*��p�H�C����[K�_a��N�+�r��N�mr$)�]W!9{�����M P���C��t�o�%� '�ܿ��:�c����]�c���0���X��+�n�C�o,'j���.�-�j���KyZt��/di��	�JdsK���8��㋹{�P>������u�ᮐ�ҵ���pse���s��ݣ�Kp�wԺ��rʳ�q���֬O� ����J mW2��Z�	Eo��7N.t�K�P��R�~��`$�~��a��0$eI[kϒI�"%�4`�VϦHǼ���x��J!��}���-	�8��	}�Q��e��-+��&� C�n�G�G��OP��&�p��te��%Uv���	��ѡNL�p�Z�"	�t��l����.��$��'�qϸ�̵Q��Y���]ʑ )@���;	F�X�c�!��2��zM�f�̯�������R��Geh���Eط����PAE��n�8�A�I�.ٲ�y#��p����=yuf[&��Ug���|8b�xT�oQ�{4r�_so���������5.C�憤�$ *+A~F������H�AEQ��H�Ā]��g��<���� %����6���B��%<k5���>�pC��PykSEYޢ����㦕��@V@�^����g�0Q7���ç��v�������i⩊�N� �j����P���+p��4�#��/QyП�<�V*��swy#̺����}�s�\��D���c$&0&Ү3}W����Cڣ��}�k'];���\_;�;�E�ܓ&��GR�Ö(PU{�:���[y|��5�]#�x�����Si��u �E�W�D�X�����|6�n��;�mD��A�K�c��B,�g�ntEY:!_�+M|�~����EvH�=��ճ�&��6<|m���������!׽ޑmC�z�"g����7A�"���b�<���)c��o��wޗv�W?���&� H��Ү��G�B���v�՟j�U~s�	{���%][w~K�����_����g0U9�wj��k�LCr�R�����-�Z*��no݂�N��0�[�_���jJ�s�`툅I���V�&�mw�j����ϟ}����;Z��g����{"��/h��D��#T�C��95���Q�M�ԑ��G2�q��4�BI�}^/��"z?W����u`��J�����53�E�Ϙ�5��)|s�n
�d��?��A�����N:����X���ÂC�+zq��N�6���X�4/��SFG����uh�}�!۲�=�EՆ�^�9�*���� �%�>>�D|������,���A��s�2�C"	J��U���̓~�	RP�����ľ�:��zkZ7p�{u���_RG4��\����fi���(��I~&�OmO�� �Uq&��5Z,po��V@uȚ�� �e�Q8t�e�&��m0��K9ʓ���l��vD�5d)ӳU^���"����eM�H!��b*xLaYI��;C��j/�qe����?F�WG�yޔ>TU#�J������8�̻����?[Eo��}Uy�9�M�A�֜+���D�{�����Vp�D?����a��o[zr���g�Q��=d1yrcȲ�Д�9����&��4}tiXbʙluCܻ�粂��.tC\�#>	;Hr�v�u�)�/1�����x�L�6��@獪�0��zR�A�%7�z0�L�?�$��l��(�e��.v���:��H�@���ښ����%�K�n�L��߶X|��BFd�"9(�6~Fn�zb��jc̣�-�
x7
�k��}�"u���2�Y� `B.͈9�Ca�	nf=�Hb�31��N��1�YJ�|��Ђ���ӰT@�1BZ�Ч3@4��ŵ]�-��
�D���Ǎ�O�kiweؠ���8f�zLa���G�[� n�o3��/��vc�~��?�o����Yo[Ć�h�|������zE�K�5��C"��j8l.�wRo��Dv�G��mL��<J�A0b<~�#v#�}����z�*X%M��E5�;�6w ��e��t)�:B��;����+5#��Dg;�8��v/f��q<�=
�t�B��	�Ӛq�V��q?���D�+�v��>�!�r�jW����(y o�:Q�N%��1~->׺Y��rS�O�.�!9+X�S�S_kfEV��)B�e�Аop񙞊�LǦtr��:���:d��if���YI}?ߘ��f�y.ZIֶD�{��r�b ��CC��΀�s(�쭚�F]r'�~o,ʹ��Ԙ�`p�LL��%&fE�K�Ӽ�]b3e��N(�Ч0�U�� /î�Gך<�)1@��D�{d��L���� �~�D���`~JV2(m��
�������xަSaZ�y���v�eC�y�)6�k�Re��k�3=CѬ��ko��Ɓ�����p%�2e�X6S#�=p� =2�Q'�D�~�L��xx��ԍH±^���Dv�]�	ht�ʑ`0�x��*���%�Gu���]Л������g>uy-��p�s� 9���O��ۤ�>M��mw��D���f��*t��|��0og;89r$h!��I��]O״�W�0ʎ��鍂2������g����_��&cn2��#>�1�)�M��e[mwC���8���jȄBr'Y�z
����R���-Ҕ�����M��;�bb���x	A �/����i��K�"��-�lo|�⨍���;�;�2��MB��N�@m{�z�̔��o��v���~�fغ1��k�+-�'���0������+,r�ߩC�_������>�0Ͷ���jX8�v��ϻ"�>+kҋ��nz'�o1O�c`M�C+����ŷ��SZS��HϜ~]r��S~�����9�OԱ�~9�~�V���O���b�����l��@���W�;�,� r!l�	o���WU��hW�3���|5Rէ���s��x�Qs8a ��ue���*�E|��Ƚp��(k6p�����VY��M����u�X1�x󥆗q�uM"�k;ߐJ�G�����J޿p
l�tg6����G@�dOS��:�3b�3�9�k_3����S��z^fW�J���g�#A��8
�|ِ5�t7ƃ�/�>l���Z��`���u��L��&d�`�u`"�.w��M�����`L�'J��٫�Ϲ�V�-��=6��d�#3?����I	��+��ӃZ۫�>��ܘ��$]3�*�x�t%�s�GѭCa;ۭ��Ix�Q�*.=����W�ҽO�y�k�����k�eH��m�@�T����Q�����~�4�*��1��:��_�v�oQ۸>��b�6�.U�%!pǁH�{�k��	���~�ζ�$+j��龯&��Ӈ�C��[��C������E�|\Y�̥9Lٗ��WnQt�GD��)�,���D#� ��c��w�>떹2#퓟��,d/\��ySآj��Q��X�)t�������V���9Z�0���v�:b|R�Q;g��n�xioTC/[���B�}=�pJ�_�y�[v|�;�]e|Ӥm#4���Z��l*�=���
�'����̜�] ��<�l�wn'8�nؙ�ӝa�R��c�xS�!���j�П��.���P2�p���?B;8���y�l�&�'�8�\O�%�<�!�3mP7�6����G��;��;!ݢ"��k��H/Zo�p�E��t�D��( �Y�mfK'�; 1>�������sX�tR�l�@>7b9����p�%�u�g��' ��s���g쳻�����x��J��9��4h_˧j ��f"e.r��p~������\2�c�,0�t�az�x��8�^V���)��,�
�Y5�ƫ��
�x�aR��<��'F��fB�V, �d%�i -\����ӫ���{�
WǠ���#���A<$���n8�ɧ�&7m���D�^E�glV'�=b�2J�<&���)���H�'�LnNT�}��exrd+jK��/�"e`��	�Ѕ
ƓvX�ɑߛ����]'de[��"�2��4�tO���{]���}?^�]7��I0�왭���c�e�U��-ɪųH*-W�+T9��p��^�ҷmt9=DݪQ@�Հz��ko-ʃ��f!�E�!-*Z�to�.쬘�e�{�����D��/���d�~y���������a������p�S�cjF�"L�V�W�z��	Ј�ڐ{:��S
�"v�	WA�L|1�'�_�3�ΐ/��Y��jQ���f��;�#!Դ#̙uLX�f��I3��%,�&��������!��i�w��GlXu{V�d�KP0TN`3Q�w2ʥʴ��d+́�)�2�H���]�x|=;�j����Rq�4"$�
/h�1�P M���3���p�i?�f��ב(����ǰ��	�0�����rvK�K�R�o�ϧIǨ��<�~됷 E���;��­��m�UOԺ�Tb?�_��R�os^�R�<�� �fv�%v>�����>��I�aپ|l��{>��||� |�|G?�z&�fL��߱�-.�P��,�(/I�T�^�`D(��$в�W�4�cu����va=��k��v��Q�lP�9�'�B��s�^��:>���:F�V��fM$=n7-4wmK�~�l�� ���wu�
ݕ���x̼���!�Sy�>�}�# E�vk��k��� ;A���{�R�]1�PI���L-0iٷ~|X?�30��߁�p��s����Q:�^s��T��F�E� �x��㰭��ؘ��"� ��:WL�7'��(1t�,��Ji��e���x" �Ȑ毰` M{���DU�h������=b��jHPY�]3a6���*#������2�`!�u���<�� λ|�)�/6>��s��~���UVVVJ�£�L�B����onӽ���	l/&	�f�o������=p�3����HF�Z��MM�LH���\��F��
u�E��q�K@ª�x�'��^����u`bX^JA�TR��O8RA�V:{�<���27�%-Fw�`1S��R��V�,�RkΧ3��C��xjY41>5����B�z��ޣK��ٻ��Tj>Լ���8��"AHܔ����a�,:��W����B9��-���KDld]Ӟ���Ӊ�`���|��:;՟����6�?f��w����y��fb� M[��n�rG��v%���wG����u��sY���k3��D�g��c�ʠ��z�4���9���"��&���*zX���@�ţ�u!�8��k�����e�,��IX&��7ד5d�@Pó ;�����|e����d��兲�%�#^����j;y�o�[���Ν�:�C���ST�X�~�S��?	���X�.�`�Zoa��B���!�c�h�q|��}6�ھ{�=H�q"L��Z�E�1Tg}�MnƳx�)��ƛ���o�y��P��G��G&+�I��a�ct	���a���+3+�V��Ð���E��w�hy⠧w���({-!n��_�aG�.#voa�,f�%�:d�(i��s3�b/MQ����~��<uG�U),� D�����2e�:k?G��iw�8l��ہ s���hp���ϴu�3=�O���E��/�5�l4|Ў��]܊�W^�뙚�{|<�_eؑ����Y9/�e�`
��#e�d����cug�HP�(�4��D#�>g�P��|�y�-W�@%�RꜟD��I�^�dR-��/U��2��.b��Q�\�d�gl&���0��E�}��V�t��uL�D.�GA�+a5����u��1���o�:y��f����E�"s��6�{�v�C�A�u���&?�%�ɳ������Ӎ��׀��fn���12�3v6��ǝvF8u�����o�-Q�ۭm��q��X�.�64,m,���meGҪ��xy�r0ߝ�J!�#��`_����p%O��n��n5�Q�F�ValE2[�Db,(���R����QZ���st�#Vch���F��/��pZ�B+�ql5bO�IS���8*�`>*@�e=�ּ]V�A�i:v����v\_D�<F��AL�0�d��'M\��8P���N��=��ݨ5�k��gظ�L��k�$j]H�̨�.��[������l�?�T#j�=�2��?��u貘�e+z=W�^L�4��s��\��+ȧ�t�]J��Ɛͷ9����b���bc(��NII�OU����b��"NCC?Q(AXpF�ƴ�F�R|ׯ�XN.�2�0�[�|-w�'�0�V�bx��<|F��`9�1~cV.5n���0J��`{�)��	 �X�z����W�.�.�R����RW�6=�0u�D�j.]E1��捳
T_������5�۳_,#�α.݄�u��F*m�H�I�Q>s���0��^�k=;�u�U'�ە%�'M>bW�9�����?g�����>Q1O,ބk'�����5B9vcK.��  ����@Mt��7.�O�:C�DAR[�(�T��Z�66-�������;NZ?���ȵh���ɋ���}d�U\Ֆ�ֆ���_rc�Eg���W�KP���d��XZ/�o}~���P��`(G=Ƌ��%<"�.����R1�FK�K��/Z��.u�]4���ɝ��&$Ls���
�ޟ ���x�堑W\ku_��l���6AM݋oZ���I+�r��3e���ߖ���{0�j}X���B�����Q�����o'����e�c�mL0Vz�{�'Fw��5��u�#�w{�>�Ѝ�[=>�8Y�]�u;��=�xj�h�.�?��oOݍ'��/Cj=�ppu�|��)�{� *�k�v������7#��^�$�.l7�2�*W��d�O�v���20Nr�1� J�Œ;e\�ww�Y*�#����v�k�bO��o;_�kO*R��W�%�1�\Vg�1�Z��c�Iu+�kZ�y�]�k���"�O���]ɐ�MH ;��W?g�6�ή��0���O�PKb��$�����l��Adb��u�W����S�Ce��K#���$��8��X+���$t/��5��4�`P��Qc ����)\�IdN���s�NL��QP��ԽeJ�k^�W�@��X�np�~����D�!�{��d5eŞ�}��������>��O��e��xy��Z�U�|~W�qw�$�yO��?�S�Zϛ!0mf����Em�%�w����Ё%�� ����D]�,]U����m� L�XJI�X��$ۅ��9!Q�����h�7U��`u������Z���3�Vlp���J��m`T�ч��F�3zU���Q�+n����������G��b���>A&`��Hȷa�JfNTD ���@\��0���# �dV�Q��>>�#�� Y�{��μ�a����VDߩ�
�4;8���1v�V��:��b4�Tn�Tx���DD#/J r�&�J��>�q�7o��7�d����<��^g�
n�b����xBp�PLU��$�{��ܺ�����ƏF�W��=|굖�<w\�:�#�7���'�V����k��:���,��V{���a���Ha��]�?�2���뺥8w���.�)�8�]����Cq(Ŋ{p(n���]>����푿{����N��;��yz������8RǨ	�m� L�eC���ï
kD���;[~�w;hU--�g��ӕ|��C��+%i��&%ΠYXX�#�G�i�{$uU"� ՝�9V���?���1<�<ڿ���=��]Gu���>n�
���z�z�:CR�k������6On�w�� WK�ZN�����U�_һT\�R@-������E�p�rr�(��V�^���@����kO'��:�&�G�]���t��-6�]>N*���-��\8)��q82��<M��0�~�	ǐ u��.ŰE�㰥���r��.��Z�/��f��gc��?׊��7:=��K�0�y{z������aFb�_���i�F�����tk�����Tɤ0���Ɇ:�o2���w,����ON�М�C.�7,����7 ��$}9,:�!��֟�^�RT~IE�p!����b�J9�T����l&�-2�,X�$�NS�&�"�5����_��oڵ� �Uz�R!��*��ߓ��6�͘��H+�R�J�#���&aI�L�k����`O��X%_�8��hj�����v��<��c�;�J��d�1͡j�_�~X�TK�R���̪~x�Cc��;�\"�
L��}��}�b�qu�4̓g�K,M��1c#?��_ڵ�a������"�8�NNV�	�����kR�qz�í�f�{J��.���ۏ�a�5+� �"�����{q�f�K�ٝs��ㄨԃb���R��mM�����0���]��O�������h���J�ZT���yeF��8�y8����\��.j7#rh���ÏrI͝\��r�v��ӵ��N�[�'r��U���J؜�����z����y�jʏ#U-��(c���t�LR	�\����x�,\/�6*�9��,p)aey���P�-ҵ� ��޾��Kri���$���~(y�b^W��:Z**�=dG�?��{,���[p�'��|��ɓ|�T�0sYBɀ��ĕj�.T���Y>]�z 2��`ܱ��]��尷�8�߿E'#A�|[f��\n�Y�
0q�nˀ>�^�n�׿�/g"�"�P����\���g����b6�P�E�yF~�'�pn��N�("�S,%-�� �xF���=��$�t��|��2�o������I�2^l�
��h���b�D������Ж
�Ͽ�oy�O�D^�>i���2>_�o�F�$Ô��n���u����߽�~?���[C_��G{[N���:��VRR���g5G9<6BWM�a��� �ǚ����J�Qÿ������"�~7�D OOH�v=�ܦ���ށ��OC�ёo��Aa�)]5�VK8*�w��p����U�7�9Ҳ�(�e���3��S?�Iu��6�;6���k��2���n4[6��k�P����C����OL�� _Z��r��`������v K�]���#7�3/���:X��׈�T	3�*F+�o('��;j�*a��}T�����}�(.R�U�����$gwOl﷮�k����!���݈ـe�hǋi�Y��h�sr�=���eڿǭ�B���,(e��!��Ͳ=&��<"F;�i㒃�#_d*W$Ũ�0�����8���l�,��ecC2a���U�[D��1E�%-3�I3˒����/8���%���:h�-Ɇ�(�iP`ڮT��3n���)�w�sf���#4�9�_�l�|����:��-��;��?� %�vG����ZO����L�K+�$$���+�y9Iz�Y���`�r՘�7W�Sr��+��C�n�R'*��">ˁ���r�z�����Ԟ��<�S���`�,:��σ��Wc��KB�`��U<��z�)���|�1N/��!�&���.�仚���4��>M5sk�vVeZ�f�齔]�`K؉�~��
�!�Ow'�Hd����5�#��̤�� e��k=<l�z��}r���>�V�ã�����VYB�썬]a��{!�ᝡ����]'��S��*R[el(S�]�/q����@��ȃ�]�(�H&�$_�o֏���/��L'Ƈ��5TA_��z�ĸي3���ͭcK�d�3lǯ@�*x]�R�Ml�FT�i�B���s��4�pY���
�N��:��°�-|@���w�M�F�6��0����n� �Q$Y2��9*�c &����o���}�=��4o��jh��Pk��5yq�)��S�� ,Uz��%[�Z�:<T�+�&mwH�
[1}�������!��p� �A�dXr�l�
?�BT���SY���4or:r�!�{[����b5���@G�@�Stf�ix�6��\4�:��g�N"NU�J;(U��է�D��R*�@��NO�[X����K�~�! ���w� E���n[��T�%�UiQ��� ��8��U���S��X�p7c���j\\8QE  y0��G7r�/���q�T�$|��M9J���y��'��$4ޭ��<������ҵB;g?��8s�w#��zU3��[�}xc(,�ۜ!���x��g2=���<�;�V�_%�fG����X#�=�B$C҆b?�&�zL������K�3U����E�/TW�,�-��@����Mu�^]
30��!m֡%�QM ��U�,sT���"�[�#��h�Rc*�'��Z�,�
C$�f,|ǵ�%�μ���y	��za2�#X�l��1,��^�0ڤ!3��*�*�LV\�M^���/�UA)*;㎻�I��hq}[%0ؚ!ڋb��46�G.�"��w%	�<�WR��[�����JDy�Ҥ�ᔼYs�:��W8�fd�[���1����Ζ� @{z���Q���_�>���!K$&�k�k2 �����!�x PDǡ|�,Xg��3���K���mM=��w��n���^zREYʔ�w�@��8`dF_�D��Ȝ��i՜��ᮆ��d}��̫@�n�|FG4���9:*��d�[�b������\>�r��(�"e�uN��V8������3��
�|A"j��ڭ��5���>H���J�'�����!�G�N�Oq�=�c�j�OC�[w^�!58�(�X¹����5��*����1��J�v��{2IE��y�66wN�wGbñP'�ҩdI�/h��©�=1Āb���G	��Ʒ��G���9�ꚻ��T��fXZI������ۤ�L8t��)Qrfz湸�m��!��H�Thaf�@�08=�q0X�J�5+	^B�ub���
ʰ��Q�:�}�AQ���@�Ϝ���F�}�狷s��)Zc|� �܀ƨ�~��a�*�P0[x�σ	���B��(r��!/�/���u� ���˅A鸔ϟq����k�V02`��[]�)��A^5��=¦]q�=�E Бo`;�0
R2�r�-y!�UC����/nX��(�n�748��f,�e�խ�m0��d�����9�7x�]���yξ�C/~�ߗڸ�3�ya�Q��s�<��>R���<F�~���4���{Ɵ~�`�fH D�J��9���:�_�1�g7�t�|�s��,A���Q������T�M�u��)�?�S��gb�����c�-a�8����;06���6U�5�7���j]�#�4��_a`�5��UƻK"��4;�Y'�k�XX����4��Q�9���*�IS�H��;:&��O�V}���W$+φIk�P{�����(2Ð�?�������a��ru`��G�qZ�f=�D��0��>�B��q��F�R�e���u��{�;!�W�V���;Ǖ1� Q�JGz��x��x%Vf3N�Jn�����+8{��������P�9��L���vK�81+�P&��iP�ݘn���ڐ���0�3>�����W��
K<������5�K%����\�i���4y��% �w��U��⸎��Hv��D��l��e�|�=���L���g����'rN��Hp$����}�g*oCE��_;\ ��S}�������[&<�ŧ����lx�h����ٞ�ld��2���ſ�����4>1Wc6���y��ÔH�6+p���A��̗̈�sR�����i�`RZ/E
��%�'�p-�p�yF�6,�tڅs# z5�l��k�7;��]oM�u$�=�n�{�́9W!��_�+k�I�:��Ȧ9s�&�z2��:]�Q& ���	������S�5k�E�l��7�x2�Ԑ�y@¯S��P�?w_l�u닓��U2	?O��?�I��k�1L���r�A���k�Hm^*F�a����pE�t�ǜ\��[���#��Г�D\R�����z�nE�f#8"�����Ł
��]���	\E���d�F<H�d4MF���X� hj��Y1�4���E3�+�4��@6�Œr򉴽*	XmjD59��b'>�=Ĉ�)h�8��-�S��9�\��im������V��&̨m�%ƋJ�6�0��a���'�G��*B�2���1Ȅj?�������>R�.I*r���y���T��d`���Ҧ��'�ĉ���fZZ�)ezN�%��3��*B��֣Zz ��lbq$�Ȓ���R�#GJ��nY���E=!͡�YG>⫔G�s����l��)�O(�;QB�ds��>C}�}J�	���ʴ~�;�:��4�D�I)�{c���Kb���nZ�Ŋa���,�@B��L�9RpF)e�R�Cc&.Hh�������.��K��u����@��a�� ��6�IҔec#X������	�;�"�Ú��i߸u�e�e��C
e�J�	V��oVcBJ3��|��ۜv	ք<^�!���xc���:��kk��'n��2����m������c�9��ٓ��ߓ�M�2큱I�6�8iÉ�511�� ������Cz�Np��vi��E��D�nV��|�Lt�D?�/�/D9��4�L�*�!��r�3�9��DG����M�r�)Ui��Rn9PD���.����>���{�˗�+ x	5��2(��˃$��D�B`��е�������&%�4��$d��?i����R��"���@�� �t�T��l����+�U�Т�/��Q�"[g�w� Z��mƷf�yv���x��3<�϶ ������IMM��M4��?jNX�4p�puO�B·t��_A`�'�A�k$�~Q %�]�b��^�<��1ނ��<�[.�҆i��'Ɯr�7O�`��8��ۻ���e�O�������~Vu��D��P�� �Nk��O�������)���v�_}�=����	�j&9K
9��Bu"lX6����@�B��b\� 7-U�����U�'P���-+}2��#qD���H&F��;����v*{��=���I��y�qy��pM�U��!Ǳ�=yJ�n��LP"�1X��T?k� ��,���QB=�{�%1q�����3�!���4'��9ҤA��'�![S�x��M�2�����J
/��;Q��)�k�_��l;o�J�'H��a�.]�Q�f�~]뷅bL6�~!9����2�4�-~B?����NT�T�+���-lFH�������
��³�4t��1���Μ��k��y�*)���+����)s^s�R�qHe�RH�� {�&"�)��Aۆ�˄U���8�� ����m�lh��`�#�D����I?���s���q����`���iq�wk8|;"�������m��f$�����y��?���>�Y+�ဳ�9ڇ�����*��K�|0+���_(L�Q����Ie�gV�WN�f|X���2x���t�(\6zG��e�o��R�F���P�\ќ�W�6���u#O�l�g�O��Mt��7{��x���� �Z�u�Y�{P�,���x��3����"|�n���LP�
�UWYc�T�S��z7���!�D_7�!O�/��LS@��T�Y7N?��e�f�cF���D��quJ|��O�*5�)��oE�"A�v/����c���q롥jk,U��Y7�>�}Y,�3K�v
�w������������2b�cRp����������������fŁN�u�l���V1��8b�AY��X�R��X��?��+��=��N�5�DQ=����\&��z��$vssER��A	p������Q���3�N�m�$�3�}Y�>ӑ����٘T?���	)��^���b�Y{��
r�e+��Kb5��E��k/ZмJ���ԕ��w�ǋ�E�F���s�t�ˬzj5 &-z��c�kF\�Ѿ���VA�]����ڗ�ׁ�y�&u���O:�F{׋�2:�����;���ppp��8����c�����U:���ܲsL�k*�jkTD`*����q\��6���JO�2�ۛ�����l��XY��)r�T5���Py'#JT��	T�`W�!gRqz����=�a���8�ɦ��i�c��"�h�GlW�������mJ�3�R6�7���=ND�9�$6�y����$���Jp����pH與b'� r��vSGk��#,r������e�}OV,Ѳ��mg}o`�O��汛�^�9�ɢr���fsȲO!���\�g	*ih�W;���/l/5��G��\����A��ON�\dg�Au�ɑ���[�4������S((H�6����lg/��򉒍�`0�g���Y�rY_�F�ll����2"����y F�o_��~�#t��%��D|�,$�6�/��B�$�z�Fn�H��kb�N'���O�l.�6��ħ����'&��4	A��-(�8|~0
�m�U��ÉV6���~g�wׁ>�����a�.�K���򒰸�'��P��^]V!p��Qs0cOAMq�r�N�@�)�
�M�t΃�t!l�
q��X���r�XR���
��ƙJ:,a}��?kk��%���E�Owa���.�L�9"*e��h	$���`� "���Oa���LP�GB�d]]c��.�Yb��ٚ�+��]B�K�� ��SC�� �����񯔘:}��Y>���v����B�����"t"�p�@�ĕ5�Ru���@5�ą�{�B��V�� � ���q�"�,������OǠ����ESߜBП��5�AY���U�u1�Q�l"#S3��!P`E���K�t�f�&R�f�O,��D�>�W��]�:�X�m�&��)}�TE�&�j/[�fݩC����b�*���lz]H�F����V�G�η*�T� �$�Z���6ÖP��r=��xTs�	�Ǳrn��ŤƆ	KL��T�,��/t��J�S�Ҏ\'���tb���.w��o��8���Qc��%����o���n�\���D&Ra�p��!�k>���L0;�|�wl|�St��E�h�����7͏���Z2��8 h����%�*�g��$�C�+F?�zC��ەQ-��S�*����b]�;(\ ��K/�PTuPn'��5���勝����{	���q�&\N:}!o��T�1����cX�,���ϳou�A�[g�y	�o��s������E�s�����H���V�5R�n��@�3^�<�5,v5��� vx�"��O�fz�����Ĺi��?,v#�۱t:����jIme�o����ל]��[D���3)8��^&r����`�����/Y����rߺyP��^����J%r㏓{S�4�z�WN��%��������=
#��H��Z(�b����w���#�s��GRi�vj5��ܻ�כn�E˺�S3�4�EoD����C�B	Vq��������M��f�ئ�%����4��	���׫v��Ƽ]�R�0	y�U]̜��{������Ӗ�o��Y�dU������Ŕ�VR����b�Ы�
�8�7���%�X.����Oug]�B�"�7h��E*+�N��P���֥n��=*�lާ�Y9$y5{N�f=����r�U���� �U���N��g߹U�m����V�B�F�w�>�L6>�!q9���w0+++�%:zz��JE��5#�-r?����%��������]sl�#J[�:>����S<w���Xe}[K-��(t��zh�8��&�*z6�.-��Q5��FS���$��k�z0+�����s�7s}+Ub�b���|Dn̢�4t���̾p��E�����"A��K�#�U1HS{6�SA����I�&�|����j���I��X
)�>{@���nS԰Tb][�����ooo���T@�oK.���ꗷ�A�_N�	���w,Z���`*�)=����ǻ���G��[ݗt��:	e]�h���R7?�V$�F�BqՕ��yA�����]�c�Խi�v/�U�%'>ZX��a���
i][�Ȭ����ŔUг�X����_DH
�1:j_G��m���x8<�M�~Cj���>�|�3kp<P*�9��Keg��k�y��k`R�E�͜N�B��h��5��'�.|����m�p�َ�ߣ�]4@-\��F)��w�~*��nl�pK0OM�S�EFX;;���M՚�w�!��z�3�: �ࢯp>y��Yp�122����]kX B� �ρ�f�����Y�HG�����|iA�D��~��j��6E#�� �җ:��(�E���0�zX�n6G|d�.c�嗦`_'���	��.hos�e�7ɚ��ۿ4˳�̚��R��p��}¼��i��"4=V�$[�nׁ���-;7���|���El���q^&���MZ���2(.�2��#��}f�ٱ�u��h��h�H2��������tjc�ĭ�~���m�}}��<�e\�C�5(|���ُn��`w{&
|�����!'�Z��) a,�z�Ȩ��O�a3�:t���Wl�7�WH�9��i:�����*r�_��e��i��:������!�=���ܺM��k�ŉ;i�9��Tʊ��i������a�sAXj},�z)��F�ٺ�8
o"��O����GJ�y�[�[1��v�1���dʗRG;\�Q2�-��O�je���0w�� (�����ż{j�5ǹz�g ��9���t^D������}}H_�U�t��ge��b� "A��Pj�5H���q�h�5�`�a!�W���f������a�������eC�&����c�K֞��V�>3���o:��mF���h�y������PF��k��o������y�c/���:�^���O����#�|>�v��أCc�8�5���I ��pik�e{������H����Bj�RܾA=�����I�۷p�M��W�f���T�R8{bwV�8pb]Xjk]���?��p��=�~��`��Z43R�v|S*���iJگ��#�a�u2�\e��8�]Є�Z�$c���6�ց���:��EG��< �Fd�0[��*/͸����:�~A'�@w��>�a��eu+G��3oI�V�_��/ڥ��:-�y?
��o��tO=�#�ٜJKk���|�ĭj���I^ID���^��S�
.����3����K7m>������zU^��ΏZ�a��P��a�@��~a���&ߞ?�q��X ���{R�c�>'!���,�/�t����	a�9�x��@���M����0tYYdj'N$���b�ʸ���5��ۣ�&`ұ�)�SOi�VX9Z%k��?'�����S�ԫ���q������#D�"7��y��6���R\	/W�8k����R��޵�n��V%�zI�1ʘ��V)�44��.:�*�o��N,oY�Fq�	(EZ�"�
��
-�SjIu6���V�5R:�g�� �Ո�Ï�$
�� 2�g�~����<T�Z����$Dsh���r�_��x֠�^>�	!�E�[�ϻM�憗��)���=4]��L��A\��TB:5JU�jaE�8����8kwܜ�?�45e}�ٳ���!:�%o�3��KU�3-oZ<���G�o]�C<xODKE_u�Nk��k�~g�m����x")�����SPP�#�x�k-=��u�ؿ�gad%B���ܿ�!����tX@FO]�9�V�|v�#��U�t�dZDI#��F��t4�G�n[�"�@�J��V����@B�^?c"��/瀦����^oI: �|F��B&�v*Wt\���F�9��F�za�W{{t�7G��hSO�]��%Mr���Ra��uP����Qd|u0W0<q���d�`DT������.�SI�&���L���;K����u�Q5	w!��]��`�ޠbU��j?RЄzd�˶9o%� `���V�*x�ٵ�ō��ʔS�����A��TX�f�Z�K+)�Ό�f����y��YZ*X����*Ү�oX����~�|"2rv������LZ�p�#���K�2��aQ�pd\�7��)î�G���#s%\�y	=��%T$+�I�$'kI*!h!Ce64���{<I�I�j#`����T���1�V;V峋'��Ǫ��eD8I�厂�n��.O����e��s\,���RP��Z���e��!na��D��@}A����J9��o�����F�C�0����j�Dgœu�I�uܗ�4���"�t��v����*a�L0��=5�L��N�����/͸�7�������2�O5ki����JP��GH�/+i����b��1���-��Kҋ�ץ�߇1\�Ld%b^���!��D3G��<s6\����a�zz����E��SI`Dl8/���gg�Л���;��V3�4|����v�L�C���u���GX�5�C2@&�H?�V[�eV< ��
����kUҼ2S� e3�����xc��! ��1P$�1Wc�����B���BhP/���xw���i �x�PV
w�/���R)�Aw�Z ���A���+�Z��][�b�_�i���+�39�tt�:o7$x�0aK��HD%���eN\{���%�Gt�S�����K0/i'}�*��XO?T�y;qf��Om�m��v="lH˽�+Ւ���M��l<�u����;8<�#1KGM��t�6���Nv*�xYDAr˹[�"��Ə9���oa��G�N�G�^03HIŽV��$W�����D�M!���||z�%��Cdr|\��Ϛ/�:��Ė�3H�����HV/H��>����pǮ�R��� �%���o섃�/��)�t)&���9ad-��Šco)���Ar�ߡRS���a�D$S�͛�ZFRgWJ�w_�q��2�����=�6ɮ5W���T��Ȋ�����$=���2�?qI(c60��M�ٓڈ/�'�Ё�6=Ȩ-��fnn�ú��26�ǌ�������� �:�NI�G@����{�bL2!m��&�E���!x��+8Jx�bE�L"^x��f���x��^=�s�{T�mu���+3�1�V���e���'���ʞ�ܻ2�&��:z��
j@K�>�=��b�G��➵�j�}Bxq��wg������gI��_����������`^�{#,��E6�A�`�k+y��D*~���xF��A@�QUAӠ�Z�̯D���l>�ț�� �)-L� ��bc÷��w�&=�#Qق�l�:B�%�_�ڪ:F���K]%��4l����>k�N\��Mɺ'?}�լ���o6h���&yq�����G�}���RIɅ��Wo9���J>��ꎿǧ�z~�8���0�/��|�!s�ƻ3Ń��.o�W^� 
 ��*	Eh��
���"jr�=#@�	K �3�K��h���J*8��F�)�f`螷�ܷ�1�7%"�;�>w�!����UPa�%���K��Ad�KU��ō�$V�Ȗ�E*7�H����w�̜��a��m�e����s|9Jt�l�k���*�¤�_��"�[Ja6������$I�_�����3�c=V���M3�F��-��257(7ñ,-g0��V�e�\�G��T�a���J� DLK=�z'�_mQAG9M�}���e����� ���&� �_�,�3��.񜝝��uL}}�����z���dˇ��J�G$�jA���%g���E��L�DAT2)yj�o?i�Ћ{��{?c�����r>X�1�Pg�1��K�=[�3�3�PQ�7�Pq`=��V���Z��>S��S{�K�������]�vL��"w�=�#9f̻DM�}�ɢQ��h�C*�D	7�r���k��>��;��O���b˷�I	�"�y�=x�Ž� ۟_�<���R0�_�y)J�cM�iyz�q\Qy�>Ƿ�@��6��0�BC}�X���fd�"g{F��6�rX��婸���^A�nnnuu]~�4*}}�_n��� ����v5u�ܿ�j	Ài'���0A�1�8����^��� �rU�r�͌��ю�k��O����Y���Y@�Z���6ŭ��Ƭ��{dXV�\�*���U25IR�f�q�����/�
���e�����	�j�v����O�����M�M�@���ab�	��0!��"G�{�)�����"_=�;�Y�w,_�1��~O����Ts��̉��M_��~��*����^�dF�L�+ ��\7e��z	�ir0>���>93�.�N�E@	�b }3�'nY�JAjo�Dt���u�����%�Մ��t�E����g6�׬�W�p��[<ԇ��l ��ӳ���-�!'���ZoNfF�A���:>U�L���8��,k/UI��W=YY�I�mlQp|�:�{ "z��t
�A�SH[�����'�����r��J����y�QU��X�e���N+���JP�O^��@��|	!��]�1/L�Z?�o��r)�'3M�p�W��ޜ�����*��^�I�J.p��%J�D�+�Ěˮ�[]g���Ð
��Q��e�W{w\фv���GwE�8��1�_��~�����_�������^�"�Ϥ�LP�Ԣ�$Ԙ����&j���xn���T�3W���� �`(���0��7�Z���έ����Aڜ<M�ی����8� �v�c����zp$��#,<�R�%K-��7��C���২ŏ�����}|2e��w;�#�A8]��(K=��,�	g6X���@	V]h������9��=@Dl�)�X��J��I��e��jrA^�G����%{/����@%�Cp9	\[Z[*�;�zQl��a)` �ͽ����woʊ��C���MWČ�o9}����I�Qa�p�1M���U�{���QI�LV�L�gX�W���#���@�咑G��˔+������j�gn�4�Eԉ;���rVJ�s�(6	fSe�fQ����W'�/�
�On988���kp���Ůf����Կk����+����e��c1�
�K�G�tE�[�q�'AO��i���n~�����Zj�{��Xc� g�y��Ἱ���=4R���!��G�����T�V �T�F����Ӟ��v��Nh����=���M�����k��C�c4շ��f~M���k�d]����h�)�&�E��P�.�|Q}Fs�@,�>d��I>.���O���X�l`�5�."��Ƕ����٪1���ʤ��� #���#�p�NC'�q�C%�"�Z�}�`|G1ӷ|h��-1м�����%�ۍ���Pc�P\M>+T8�rJ�,�`xP�k�iM��;�"�m��&��4^���.y�2�����`�XS%�[�~ѭ�W���`#���ȳ�Ué"t��"E�����Lj��⣅Q�q���ݒ�\�F�7�+=�:�����3����c���r�>)�w\� ��� td�T����u�h������Г�o8����2�*�����b��م�6�V�K ��ҩ-t��	��F�,���s+g�̋�G�&�<%�.�18,&�Z���Q���gƉ��&�&��N�d#��7-�a��J���
�,���ϙo)45n�rw��in4��}��[�<>9iZM�4��� �GH�+����#n�m�	]r���� zU��`�B���J�|��3'nr����'6ق��??ZJM��!�8�=8����H%���Ө��}�2*Z���]nJ7r.�w�K�M�?"��Fc�,I ��� YG�_+f����PQ;���0йv�"	3��(��� ���wZ��r������tc�)N��Vpv:���\�6��_�J��t����(v�W��w�ǳ�M��}����9�h5�f9���Zw���'�Q,�X�R͚��~���>���!�Ӗ(��e��Z2'��o�R�#0YD��Lrѧ0r/WC���:���`�N���tŤ>
�����R(��uBW瑍�g���Jٞ��%���P�5N��۸������]��-��^4ђ����aTsp��唝I�*R�*ܗAh�����s�osf����"mS��׭^��f�!kݖ-��#  �!@�uv��y׍>k�����w\�~��'{;��C�~���&�Gq�JN�N����F��)�n�V����X
�}8,��#�ֺ��[�;:�o�kkk;�r�,�����u�k��|?�� GU��a�O,ǚ�"���絧�`zo?�>��}͉µ^tM)��,{d��`0Ϣ�p�tN>��|��È��Q�"hg���_d�]��N\]�h���|��ar�f%XQGW�G NI��-�x�"�F����,����V�o��)(�t�U��t�e�]^�}�3��wĩ���@F�DA����� �9�U��;\ω�kkv�e�Kz���]��ͨ�J	RJ����Y�H˿S��y0 9�uN��!�{��m�FE��k:&n�zI�����[l��WѪ�b96���Q��H�Ɔ����b���}�s�]���$�^��Z�x�~�K�ۤ>:��Ey�eխ!-�?3ju����Bۼ�(-R�[2�¦��DoV�,4eE��[��;��	YAA���kT ��l��T�����o�xJ(�U�؂+�+���Z�,���0�&��wЗ����N�񫡭��0�v��0ps|4���w�Q�heNG@���1RX���>�9R��iEG�7�\<��I����Eh�+���t_)���Ӧ&��v�O�Y?���?@�M���`�G������8��|$ɍ���/�v�A{���ǧ.m~��r�ӹ'd%{��\�V5F��wv���y�ek �A�buN��� �b�0TC#�=6�d���	���3��������6HP�=�J��@�A�X�����1"��Mj��e2j]�T�Ɖ��]cU��Ƽ>~��?����{�Õ��L��N"��n�� ��Ӳ@� �GA`X���P�Uf���?0�f�*��Ɖb��;�e|�������C���E鲨=�Rju�<ֿUw�.�/��[|`/��,
?��<#	�U����_Ҥ���x�_O�7�����ͅ��"{ڽ1n�!���茌c�^?�>�G���8Q�|oB0Q��\�"#/��H�U��Fƃ����nk�\7t�@�4�Bj_4xn6!%��������"��!8���k�]�`c�[b���8m�jř�����(V����ώ7G`w������O�z��e2A^*�TM+ߢ�z0�������Ꮔނ���dҧ��}}�j���
j��~�,��N���f�x��a���_�C
~��g�;�bw��Vc�^B�B��JY��/��5��gY�	�b���8��c��[5��LT��S&��]m�S�aS�5L~�YS��'P-hNFF�Q-e� _�6�ښ�C��t�^M��)�T��7��Gi|�h��,=<� ƿ�j�.{����P C � mM�[dW4E��a����:�b����7�e~��9O��\@3i�e���(��P槠��[��D��i�5�F�������6�~���Ė+�'����`�ַ��(� ���u�ҪP~Tk\�o��֨]�g	��w_���ض.����(���>��V�.�NC�%$��>S���4�����"��RN�3�a�V���"{37u�����8|��1�0{7h����x���{5/��g,����h�J%N��I+�x9��i�����;��\̍���;��m�DF������i���e!��	vX�kdg����&	�SM�$D� y�����g���׿���NW�-�Ɛg�O���co�*a�
�ͽ���5�=��\^^=<��5'ڙN8_Dg�$�U�k��:��)�h��Y���H}����_"x�8M�=�̦w���6��2����o�+u��}r[��^�W��T�Zv���=�����p_em�4�=k���*G�:hN�YB7�E�4�f�&9���������������}ތ�֟������7�L�"����.�>����2ǳ�f������i]W�X��B�|���y������@�=u#9!��+�(;�[G�:��ae؟#������Y[
��aT�!������/�V�h^1s���	� z�`AD�:�u!��?%�<�e@��ֆ_�)��$��D����n���AJ��i��F�;��;�=�c���Yk�����a��F�],�9f��M6j�n�)+$$̂:IV�&�����0a#�ǣ�����]p=*+ac�+��;A���5F6���-ʤ@�6��s��zq��ϳI椝���m�1k�I��>��JDp�b�P��н���C�2��}¢�/�0���u99v�=�B�e�u��l ���H�����pݰ��&�/n�WS�v<��ޫ�!,q�Bu����	u;o��X�K�����?j�rh��%	N?�8T��L����W-��7��M�EHX���ձ����@�O7���Ѱ����l���1�������Ht�)�2��C��+�$�B�rv:�a�&�<��|�+����S�t�;0����v�9���������r�Z�}-���Q��n6݌��BQ�P�jZ�K$�O�I'/�9p�?��d<U
{wԚ� *�o��x��"�4�+����wiL�⅒�n��,,�M=*�˩;�U��J��4�'���mxk4���xƮ��׷�n@h�KJEw(ʺ�V:�=&L�ĒSWю�a&&>�Ѷ������&��~���}���2�u�lN*��4ˠ���n�)J�����i�˓E{0��|�>��+�A��D�~��܍ݫ�J�y"a���`p
�2�8�(߯C!Hy���)5I�%�%�HN����"/'>"���ގ�P�+�g�r�]lpd������+��!4+�q 4z������>�JB��|��QBP7��v���u>����sؽ�^�J����On\�8Øߥ���<�������MR&�a�dAk��@�$mKhrՏ�vj`�f��?�
�I��Jx��I%�+��t�W���s�.�U�����G��x�r�T��2��8�h�8��J��"X*��Q׫,%�o�ii�-ܰ��U�7V ^���{7�#-�����GZճ58)E1Er`}����_�idNv�t�?/r�׉�eޛ�o�u�|��N1��q!�K?�|��T@)��37:2R�^�Lۮ��h]��`���F�y8�_p8
Y��u.P:E��5*�R
r4\⚢��j��V���41BR�"3�T�}ENFcg���D�8.s�]�����b�+��O���I$�q|a��I�B�0<єG	��o_T,ٳ4����h�zP �2�|�����ZR��i�R=�1�cd$5C���	G�"^S �/@|9��O�<jI�;{�l�o�s�Q�1�)\<t��h�{�c�!�2�U��t��Z�M1L��^dف�Z���p��Km�Ä/�ܺ"��-ܝ��WǞ���>aə�s�*�Z��(!'o}
j������S����KP�7d���e��s��5�0:��B#m�����7��}�a�ѭ&ۜ-�|��}�ұA������/��qښ02ΦK���;�7A������}����;��^,n����6�+>ʨ�T���@���]\�+R0�C_\ɗ�}��4mt�t =3rp��E�7�9��3v��n��0��6Dp`���졖�K��>��c�*!���>�"������-�f�U���H�n)�
�>���<��`@ �:�B}EߠG���'���mx` ��ؓ6wg��Q)�z�᫬�:����|��?ˤs9�b�>
4N��.�=^R����?}^���c1�\'pv~ҳtZ/�E��bAI��7(@U΀@˳Q��i�����F_k�烷FE�"R^QP�h�>gJ���������񾟱���I�"4�bBOe2u@P��\#�f$�U3Yk����1��[§����P�4��8�ś��?n�"�r�
�9�?��k���S�0��'�x@}���M�:������LC�T�}R_���A�J��{�D��J����d�#�G~��˿4}���YG$_��ۙb��QY�N�]*I���@�j��z�G�Vc�Ha���'N:{��C������0�B��I?C=��@�~O�c*eE��
�`ӕ2�ЮqW�����PW8[�a�����=ܦj��2!�u�(���</U�m\Dl�WN�����8�$���N�y/�<N�U�c���F�:�<���!�شȠ�Ǝ�w���j#��^ֻ��;���1�q:tΌFySWE��h=��A���������
@��� s�������<�(_�,�87����嫀ۇZ<�p:�>�W�=�}���8Ѧ���ԕ�(SY��|1-���dc��9�Ͼ�H�0���>\dN񛶬Q/V��ޟ�v��r���e(��[g��Ag�nA��;&��#wT��z�Am�_���Y99C��9��vچ:�@��vB�:�I:�D%�I�CO�����W��o;���y��dՁ�Ӷ��}%�-SA��u���wݫ�0�NH�Ъ�D�Z�Sw2l�	�]����Ң\6�l�\����(}�}�I����S��d��?�ocz5b�����L�U$,Z�����mʭ����M��Y%ӡ�2!�9.w|q5Rk���w���8:K�C=��Cե����8�䉒O��Tq"���5v���Ǡ���td�@�n�7
g6�Y�)�V����[b�����ar�#�S�ݒ�~�s\D��Cq_U:A �3��#Sg��n��[2���J����w:��.�U���I�4R�cq�R�䞍��i6Z��a�`��y+���r-��p ��N�.W[�l���+ld!u���Ю��t��֐I�'G�ث=����T�#0 &�Z6/xf��Ex���T՟{M�����̪ta41t�@[�xyE��B��>�`/��wY~��N{M���NY	�͑��"�D-��B(�Q�aЩ�4��+l]RC�S�8=T�H⸪H���d�4$�Yb���X�I�"��}_���l.~o[WZ{`�c���.V�8<�畜c��k�㘄2�&+&r�M�����f[�i��R�ᤀQ
_�J>jz��� ~{������u��
���v;�~U2(�@bzu#~ж�d0�]���|+�rÖ��U����D�A�k��ń�)Kmm���F7������S�We��cp�F����h����+NpE�e�k��=WOrӭ��VȨ[�hL['��lN�U�v^XfG�=5^4k��뱙��b�V�tܮ6�����I	=a�p�E�E+_��ג�N����]1����\ཽ�"�'e*������Ɩo1�|Mf�}D�w�J��,�sYVDP��4,��@9� ���2��"����:�04��`b�]qh��t�~�=�q���֢kA���h�on����j�U�>�Y���084*��u��1
q~����{�=18���VhB�~�x�^}�D��/��F�~���A���/Q�M��օFu��k�"��!�/��*�颁��;�eL�o��"�L�I��>�+�����,t�z�P=r��?�_r��<-H���ȟ�H�1�G�w]�؈uw��{�9R)���r� {J����ˠ�D�{w����ǣ��B=G7.�q{Bc��9�|��E]��WBI���:<ѿJt�Re:��Agq?�?��SC�阢|vn��+k(�nRm��?n�yy�NvHx�(��DB��4� �cos)��u�y�d��[�O-+T�5�t��.Z1�$З�,^��M$��E�;�%q�7I�,s���_�����G� %�Z�j֦R�!�{HA���Z#� ����*���u���
����gFH[��'��cQ�Q�*v5HрF�|1~x3b�"܆̈�y�!�?�立���(�N�Ge���)��j�Õ�h_U���q�;�׃�M|����vv���|����d�;�ĮO7�Զ�5��0�|��Q��|�ߝ�� ߁��R�rca!P�����-/�2�A�E�%�w��
��Pv�	8C'�MH��~Ⴍ�6�`=��`6M���讓�~�x���d%�Յ�w������7'dgc�����K�Qy�K�N�u�d���������;QE���b>�T��'���P����!�0�C�\���Szĳ���)���詪���q��1���o��J�.�C��>�N|㔡C�E���I���)���,ʒo3�)bt���s�6A	�_ n�t"RbZA�2�?�S�7h`^�8�߅��_u5+x��*ΡX$Z�_$%x� ��D�����_�_wd���#XR�#,S�6���^��� ����t	'��JO��e}w�XJ'�kCG\�fI�&��so���zm�ߐKZ�q� 8cߍ��Hs' Ţx�k<��jU����	����4��t:��_����21���(	}�,$�����E�5z�X�J$?�$�@��TCc�&M#4�����t�N׼6_߾������G��9%�W��$����=8���v�n����ס�Q�_�S�[h��^��;|��5��7�z��_���e~��iӌ(Y�ׂ�a���2&����x�X�OS�|��'���*y���<0>�:����N�.\�E�;�@���3>yx���w{�o�j������#m!���<o
�]��%��1�m�˱G��V�$U����������:ܲ����:��	���ϼ�?�dF�����0�>q��|�e���+�
�2��.DN
�h}e������F�J�+~�O�V���.���B�L/Q��%���ш�b&�9.�9�Ș�c�C�����+H=��4I:�L�q�,q)�;:ț��(a��	p����^�u�4��K���$$�^��;�����W#(dDG�IGNŬ�;Y�~|]�yId	��~�B��LVv��1�NF򎈚��s�)K��	�T��NO���ߠ!k�����0m�Qf#츾@{�ۨ�[3@�❠�ɦ����tu��y����5%����湛����0)�[Y�y��27��B�?�\27�obp��i�W 	ees&T޿��@��_Ԗ�t ��8ͺc������ 6[�A*��,��L$��#��`���!HDiX$\vcB�rg�R����a3���!�e�c� ����:]KRx��#x;^�Jl�M�Bd��-E��Y��Z&���/S*���P�\WE��w}��	W�����S}S��U��Q]:Aw���T7�N}�+�-_���Q�ޓ^=��2Z�C��@�?���̫f�S�wkD��P�ye�b�u@��[?��m9~w|�P
ԤI��}(x�^��-?�|�?c��l�[�mʯ��G�ut������&}�j��y̨^"(�xq�!6�.�V��~����d_�O�+�a
����c����<|��y�u[߾i�n��schTzu�Vk�
�����L��,�g
ë�Z�3x�m�����WoYgf)J���C/����Ҷ�(^� �.�E`,*s�j����A�!S���ח�/�&�,L����k��m�Ir.�g�*u
�����ԓ���ɱi�Vc;����#UEI=���� �㵆>��Ge���9��?����Φ�/��R�h�(���2����Sk�0Y���-@�j\��|zy/� �ՙ՚S����D��6��?�^�T��QjY�x]��mo��SϦN��rԣ_�_q8]$��``�"��oN6���/��Kҫ��f�ݦ�鍨��8����Cǔ m�ы�߫��;�T��$s6T�ᬾ¦|xM���Av*��b>Ui��}�/\vp�A%�{���xB���H��ZL�°��֌�;�D�PR�@���k��A|i�W���@{'W$.���d�u~�|q�O�t����p�ߎ���Þh�;�ku�輪~�$<ڇ�S��4�t.Otg��9C�hɻ_�P�����.d����m�¯��Rp��=Z�����q�G����a.��8���PC��R�[:��w߫�\��v��N��8�cᏑA߻�;���$��2����ﵵ���,���t�|���E,�$�x!��z�zW��Y>q�ktt��Hw�P�z���1�����=0�!ܨ��6"?+J��*�����F��I� �1	)��Y��N�����
L����Vکw�]���#�!_l�úM�� )ti�e"���SÙ�5�E�$:eaS�B��fN���n%��^
m�W�:�5߁�e `" �O��r�w�$��
�%�v�9SIҪ�ز�G�ך3B'����þ�ـ�뽜�{��*tZ�LW`ZQ]��h�v �}�$�W[.��fHW�c4��\�����RV;n�j���r���s���uU���Q)X���.P*-WJH\~�.5f}����ax�M�<o�,�:�7�.hEj��]�ARq!1kQ�6qqj�a�)2��D�1
ĻǾ�ߡ�
	����s�oQP�=zn��cIqP�t�� Sn�m&����1���C ��4K�b
2+2�_��:�#����T�����<��n$��u��:&�dx�����(Uq��6I�a�(aB�uM7�rO�ĽW����0wzҟ������ߖ'N4~�#1yF�3g忑�{��I�h�f�ONk����1><E�(fM���Rb�_x��� �6s>~�}�+�K��X෎!��q'ѧu��"��������s�0 +l�W��{�ܑѱ��kظV��6wx�� �I�����}���|*���SGM�%gl⋆��~�(7������	�Fބ�
�63d�:�'�k*
������2i:k���v�#�k���>O���1�ll�]{׊�Ѷ�fK�%�wv<b?�*���(�q����%��s��xG������${�w8�a�n_�C�./&��}��2H�:��%�#n�C���U��ޓ���զ����=�S�q�Ĺ�.�. ���TF��xIp�K�W'���7[�f�e�_�,+����1��!,������{�S�@"4��-�e$��<�c@"
)����r0֍HcS���Us�R�t!�E��T��n�� a!����7;��3>�c�؊D��>�nF|3���J��y�Go�L�p@��r������ۊCR-������f���E�ۉCSE�|�=~ ��$C@�'���R���qw�6�/�y:�Hֽӿ�Ee����Ns1�)D В���qv��&�wa"OS����>�Ɉ�åٟ��%q1��C�,�X#3Zm}������z�8� �塺�c��1{]���^��:������g�����߲�.���X�y�2{n�����{�ƣ}{�2z��c�����4tf�Q�cc0>II��gj���H����#F�<��$����I�7��4Z��#"kJ%-5j�M��u�(�LY��ܟ��F/���|L�9�n������DI������-xߞ;��[�T��Q����t[���<��0�R;�*]�����J�vU���|E,tԪ>��o�B_��7{�E%Cq��5r� ?֒8F����q&�}ϯ�y�s�\G��o�����SvDVD"�Ӷf3>|؍��œe�ŝ�p�H��e��S	r"ʕ�m!�о��P���Cl�p����<3E1�(�i��@Ey�p���KP� �S����6��
@�@���4 
�f
���jOX�wT[ɭ�9�F����jI�@},1n�:DrV��'|��ϗ�ǀ¿"�v�b+�~��kݸ ��㔥2׮�][�2�������`�q���_u-j�܌3>���'���Gu��S�Q���[	,T_��>��VfĠ���]~�]�����s���c�NSz���ڥ% n6y6!W�#�,FApu���>H� j�K�cG�'bc��2}���Z#3שd��u�SB����IH���2�:�*h�Ӡ�$�7q�H�uU��VL	p��%�ori�(i}�R�J+I9�H @/r�����c�v���J^��x�,U��d�H����r�D�E�̗�`k��m؉[��o��������9�aX�@g��;��'�Kr�)�s�c�9���ט���>�"��e��^��<�Jؘ��RH�)v�;
����~���ƫO�C�b���y=�8L]]_K4�4�!m�<��}�;Fcq2%x�FZ{x��a�>qr�������}K����c}����#q��A^�%�*��49+u�4�G�f���n��9�fF<���WsZ��=���m:��os��y�֖~����`Z,�m!�b9��ӳ��
����R�=^+$$e$�?��ga(p���N"�b��`��fK�����P��	C�bҫY|��H�
�?����w�s�����	� >]�ՎkP���u��3a|���Tnl����M�լ�q�wR�f�Ιj�R�y�9T������8s��{X!�֮���m�ݶ�Ñ ����x��=Uu}w��`��)
��gpʾ���]e���
����{���l��	�x1�[khǖi8e��^�fd�X͚Dt�J�3�\0�q���FƝ�ᡚ��L����\���<��e����ycc�՘z���	!#P�x(�#e��4���X�:8�J5P~�T�z!#	#琐��!�=d]*��!֋U���}�zC�zY��e6���3v�i)9:�.r�)��lk�^�r2j���}'(C�b�;C���NS�C[��!<%��������]sI#��D݆k�=6N>�/z�hCk�ɥJ�4}�uߧ��F�Y�u� �z�����D�Q
=��'�&������s'_z�g���W����E+~��!XE7�|���A��X	$�m|π��x��i�%]�-|�*�����%ԮD�u�ׁF퓤Ү���m��Z>ue�)^>v|���f�V�k�
�R���
y.�8��ad�X�Re��!s "�u���,4N�~O_����o����DD�q�Wr����hf�)欽�o�u���zo����>iZ߉���De/O!��c�}��b��f�TY;E����5�68޼*)��UD���A���Ƞ�7�tn�{�wOwf�'��9Qׅ�6���~x����u뗝��1?U�מw��0�ӘՓ��.�������盺�4���r�����c�S�a8��7�IS�iIڦ����,�����vVs�I�!���q䃵`����ڳ3ǀP׌��m��,��͡e][��'4�d_<%�B��mǤ����z�Ja����H�)���oO��w���`Ɉ��b�c��D��v��#�u���9��vd�x�F�߇�)8�L���}d#�L@L�Y�r�lL�!�Ͽ�s�(�O��nwM��(���_#Z�(���8^�0���!��S������:{���:Kgl�[H�U�W7jڏL�� XhP�-^���ɻ\-Ւ���Nc*�ҥ �D����Υ�<�c����aSm`�p�����9� -�Y_.\�yrs�lO�5}z��aq��BL�ar��r�q ac��F��8�M�*>XI�3sc�B>J��~����x�9�{]�.LZ���Q�XBQz@��O�3��B, ��e��o�ԭ]a+��_�?���>���^��3I�~���12�&^�q8���~5�vZ��P�{���7Q���h9�<����?����~<t�����:�x�1�v��M�@���q�#���:�Ă�����_%G�ίiP�˜R��R�j��7���-�aj���:���PX��%H� �"OhmE��ʋ�/�]��Yk��A[��H���FC4R���R>t�+� ����7cx�5"Y���s8�ߠ��9\�Cq�o��4�2�0_��k�Դl�V��դ t�j��� ��5A�����Waxc���q|��:*��o��w�����Bɘ�N�����C�҈f`e�����.}�h�ؖ���&,{vI��0:���fԗ�˟:�����{���2����~�0f�<���	J}�n��M�cr��o������kU��kWXf6��d��,��7]5����i������oU�_%��C�Ʃ�q� �W�p��;�M���M��s<������~-\�MKS��S�֊&��.�;#�Q�W�DE���g����z��|��}�cF�LR?6��e�A7����wq\�&?w�F6�hS����LC��RA�GYI���N���(E54!��e��uVߎ�v�����A�7�#���#��[σLjx?i��oq!n;��aI.���WL�����É���G��b�5�5O'���ҫ���̗�NaX;���
]�5�uě��~�dc�ȖA'B��m8�!�E�Օ/����k��Ê�L�X�&g��U��&�\V���Q��(b)b%���eBӾ4u}�S�\��_�l
����.�i�9����L���^�o��D1NX,6قW6�Q�y��w���s`���1!��]c���LyQ��i��2ȓ�� ���6�V﹖7���_&�'��{K�'ǲ�b	��V-�*�����W��p��۸ZZ�x�l�{�BF1��b��6���[^Si��w0��9�����J�.��b{�r�|���K�Y��<i�2XhCPh��*[�Թ�I��as:5�j�y"���QQ[���$�z?{/�<}zX������M�DT�||�Vz�X4����8)z�k����a�V����x�?��v�O�8�:6Ƥ�w�Uv��U��p8��%��+��N�z��_�����e� ƕ8�/F@���D\c�w~�9)Ș���$�u���y
	�d�[p��or�T��d�l.t�56W��wpWs���D�2Ml���@�ʨ��jhY3Cc``�Z:�v�]�`�;펠'	['TW&���q??k`��$��69��̃�H��~�3��g�UÑe�nU��R�ؑ`�m�7�X�c�S�9�I6s��򵄔e'�Rx�,+�)gt�r�[��Y��o'ʏ&�WY>��t+W��N�^�xG�(��_�B�yknMb��y;��W���m4�	����up�N�[F����϶�����+��ovW�v^�v͝��<=~�	�w�i���@�.��<��\<HwL�w�����$����7��=U�->u^��^��Y��ikǦ!U�g]A��֩�hZOV�ޚ��*\�khk�����AOu��~�L�t����|.F�T�r<����.ܵ�V�&#��% �j���6��w��(�	���fy��411�;C��k�"q}���G�va� ٤�_z�fCb��i.�V�>w�`��
	CT���.��ʿ�]?Ef��pc��,rТ��"V���-:m�lŔ5�����U)@�#M���.��7�9�:�ꕳ^�S�������
U9TM�_�����6���	���B����R\�9�y���)@P�<6ˀw����Ab��
6<)�ȺxS�J{�eN;���Ǆq�Ee>}�o�S� �c/�E;��3�Z�(�\�����	�ͤ���>loe����tݠXlo+*п���;,���Ț`1���9��\�
�ߖ�m�&�����ԡ�i�nqZ�VU���_��	ˮ�7y��3vKe��-Y�G�v]�JZ�b~�ѵ0�JaJ��-�ϲK�Hl5F�4ٿ��E_���������#pDC���L1�] �=j#+[+G�Fn�LQ9��$�N'��B�>x9	^+�2k]/rp�t��������i�@![O��U�4Y7���x���k[�l#B���s�贊)��֟ �"�+�a�g�s����C��]�z���5����~�D���%�����ӑ��7no�e.���3IO%�������N�ݰp��t���S�+�G�#E'BʻՖ�U���T(=Ρ�]u4y��ETr�R��H����'�Z��#�F�*c�-J���<��/v1����L	K�\-���|"j�Xg�7��%)��[�zƏ$��$��p�Z��~�=���1�7�w�V���/ٵ�-�7?�{h�ix]��|=�� Lp^�߽&��
k�n+��;���N��yh��:m�j�L�[�c�K1�mȝ~d��5�3��-w6
X�W��uB�<�������'C3�����-U9�|�h����"@-�B"�w���M����QR"?���~�Hkb�n-�Ū��lC ,$kQ6�Z��Te��J����6j�AT����7�I�3��^;�H����j���ȴw���'�u�p�Ҷh�Y	��3+����߬g��oz��7�dK����,�y��������,�<����Ǫ��r'a���+q��s���7�����G���i����z�V2:����Q8h��%� ��:��R7�3�!�Ɨ�Ό��>Ը��9�-b�s���5��Uy�$U�6���Ͳm�eh�fi�vta�!��J��h2G��c��)I{���Py)n�Mn	[ߎ�I�a�9.zd�o�*�+7��zL��Ȳ���a��,����Q�Զn��hWR�xz8�kd�$O{����)�����(��,����t���x�����$M��3�8Õfv-�u���N�#�I�����������	�l\��
p�k�x�-W��D��\�C��(��Im�w�w��7��We����g�̽�;��x�h/#B_��~�T�c<����=��'�4%3��Һ��/�1�H�x���̭�p(E����w(���ȶ��P 1�����
f@F'Ū��� �V�Zj-x�V}��@zS� ���vG Xl�%�/��؛.1`3���)�y.� I�Qp{?��d`���w�>��{���M�D��o�TKJz���I0޿�ѐ|$,[4���?��Z��?��QBu<*D<�Y���ʧJu��?"܁C�OV��u����LaYg�qu�I�䬽K�x.��ԥ�+@�n��ɨ�n�R�znt���f��>Nd��J}��Rx��3�Y9}(���ɏŽ���SE�f�>���xF ����w�H5�j X���7Nn��\�H�󟲉j�3îo3Y +�$�'��7��70��]C�Ϲ���^��������o�KX�d�kRï�^�}^���C����T�{@�4�A��&{i�=�R#�4�
&;j�� ����VLa�ek�7?��K37n�Čc���=�|���RS��ݞ���M�BԈק���O�:B��s��n'����0�x�G\"έ��R�M�������� wL�UW�����"~7<����ܦk�L|�+��J�N�'��y�Uش�đ�&7��
_�� G���OI�[ߐ��^1�S�}�"�����tz>Bg��{
�ۣ�4����%��Y���o���J��c�J�l^2!�ޮ���2/t��,���ڗ��Ȱ�R&�4�@���*���]�c;9;#�蜫��]OҪ�8�o�V��&��|����%(�����v�����@/��ļ�Lx%%�m�;��� ��f�k6��WD��x��gW���[Kj�����u|*��{Ls��0�[��� ==rG�@﷕�w�"�ǲ'��#�z�LPW~J3e���n�Tm� ��Tb+T���䚝����k��@o��_Wa�*IۤJ)i�C+
�`�3K{�WP���נ0l߿�{��sg` ��2q��Sv�g�͌V�:X�����-ŊoG�I$khm��m�H��ǷT��a�$�S@�.�|��_��,#u$ymz�w��{�ȓ}���L���J~}]7���!�b(���O��F6�z��j�$�@�0D�+�gg$QoT5Ol�6�3�B_$�u/y�����������3Yn��Ͽ�1����4�OX��k%oP�Uv������'W���{C���c\d���s����*�V�+���Y��Y��\N�Y]����p�0��;�YE�����,:��[�֟&mܳrr@�QJe�{ P�g�z���}ޜJA�B ,�2d�b�ĕւ�K�֥���*���W�#�(���Z>�22�1	�z$�NO�O�k�7E�I8D�Y�1Mf�vQ`YB!��n�2u7��~�)�����K;a�N��f}}nW�+����7��&�_�e�x��Y'o��t�X���S0Bׂf�gN`��a�Ǘ��f:=˃	�B���vW@�+l�[�f2U�k������UD@~��$alj�p��D� �]�� �&}�)�w��[~9c�^�\��m�c��#ֶ�����+�/�q6QZ|0}W��+�#0�M�C���Jh�������9��� s��ht;"iil\�'�i��ۦ�-���}AZ�A�5�DAN|+�y�'�+L8��o��7!�LtD�e��%?�k#�|�rү�ŹI�����_�"�]4�Ռ������.-�p&����m�����몰 ������t�)[<S��MR��jA�k��X�I���(U�+���x�@¿�̹4Y�Ę�-��O�Wc-e�!��H�rk'(V�k�!�e�._��\�@)�QEas����Q�������jC!Ѕ���20��67wꎈ3�F��W��ٶ?VR�6��j5�:��n��W�HVrrr��r�
��ݪ~"�Otaf����*���,3���{�wگ���=��n67�n~Pd�C6����4=�ZK�#`�>1G
���<3�Z�H�z�,�GO1�@F���� �x1�U��.����W7LU�Ȓ�,VA�V�8�C�!��A�B���~�J�Z�����޾������+���ϒ�$�#X�Nk�`^�Kp��`zO�D���6l�ǒ�ۚ��K<gN�F
�?�8:���x��Q��R�c��$��/�V�����m���?uѠ�|sd���;�[��M��d�gt��oT%ŇK�v����m�f�x���u�.O�?h�)L��u�c�@K��-���W�.g�JR&�YG4�J���'�]���"NiT��s��{�]��{/��GhK�4%���ND�zWG:2^�VYg����?y>���d:j~�}�������o��j��d���j�I�=]7�-��C9:G��:+[5����:�͙`��&� <�0d�F���C�]�W/��Z~VT~�I_��UK�Ƌ������A���Q���I�CHM6�ǚcX6��xUU
2�RY��d��H��V�u���\�M��D���P3�fڏ=�\a��GF�3��������׶���Fpe��p�O4/A Ў���j���\;W���#$1�{�b�8�q�%N��41	�/�6���̵l(Ңl�{ג�mLB �O�I��^��}�ڞ*�&{![;��q�����_���5�!3E���M-m�a��C�%+���h��m�)�?5��rsj�"~�N@�ZW�$�F��ճ���/"��}���@d�ͤ\g�/�<;����Ҝ�[�N�4:��yP��2�R��o~WO��S�	��ؽwڏL�j����͝�M�[N�"�W�*�R��c�j0�ii'���D��C�]��%��&�x1��#(�Bh�.*���ϒ�	���O_�������
	N���<B���_d��ڣ}�������Է/P8u<�/V�U�ˉ\�j�QUD+�s�j�0��r�Ro$�|�5�G�.�C%���˗]7��v�dF�T|ŷ�bJ��أ^*@�����UZ^S��T�a\*�\x�-���ֽ���CG�����J�nzʃ1=NC���������ӣ�6M"���'�np"��>�+����?n������ز/&����(�b�o;]���NXc[ꈓ�-@�ޢ�} �a�{;�Z��K�(Ǡ�]�\4!A.���>�詓�H���ie]�sp��/��2�|
o*��frܹ��вqI���e8(���yǌG���o��rY=�%\c�QFB�I�)5����pQ��q�0�JxU�S�YY#��vB��G�h`�돛bJX���vN�@Ͽ�5�`�zr�K�ʾ��91�d��	Jh�vw���s��a"ݾ�dh�Ѣ��2�q{�3�:�>�Ϧ m��PC{��UX蛘K'ae��ľ�wh�er�e��Ge'�tKQFeڴ��R?c=����fpJ#3@����|�+%��������G�5�7�c�xZ��e�Z����3'[����Oh��C�~m��;ee|���Q�1�YԄ@m�֮�>I��e������3Q�ߚ���$҆������9w=����ը�>Eu� /K��98�q2�XM����U9҄}��ш6}�9��O9�r�yb�'�$@���%s�����?><�SO�1��+�\=��:~�$���=c�6�����C�-`V��M����� �7O�{��HB�Q���q�2�w����e]�I��s��c���p9q1�}g�\5���s�쥱O�����!�*v�ذtB��B���>�Z�$W�zr�.�2�)k��sy|zs��Y	�i9�ö��a8��N�nfR�ܬ��y�=�x����<�������Lշ��`��aI���;�,CX�@�P�B�Z'%�.���j�w���kg6�zD>0o[gI^Gr���5�+9f!��V���@��_u�"��ow'��P��~ N�d��*ϥ;Ԅ1�orv��A��
�b-(��`�;![�^�\i�ѵbP/*��3We��b��u�QQv]�p@J:���fh�%���n�n��)�{(��n���y���˚��s��׾~{�}nZ�lPBb͞�`�{�֫�ݤ~~O������5���G��_|�_��~��D��agg7��Q�2���2��%��V�-����W�B7�2�a�F����~��~~�
A�N�+�Ȭ>�������5��﹍,\,8c�Yܭ�y�2#�[`���O0��I�Ӊ�G�1��A
�j*àpN�k.�`��?��ն_��Y���ܮֶۼ�ҔX�������Q��@��Z_4���	ER��c��TJVL�3%U����	�����@l�:��t����x��m��pT��`���(�n ��l|`�Z��-IV��������[V��7g�֣���S�ߩ6�q��
�l����� i#5�ƺם��OS.���pK��;w��r�ł6�S�ؾ ��8��;n���>�B��E��1h����C�k��R�]�IT�5��zYP�4� L�L���>8�娼J{�[dLW>5fVk�v��z���g<�o���m�����Z�ꙠvE$��:+��m��@��+=�"<�5Yz��Q�lf��y0+O˸6����h�n�����M�e���g|�Vu4���}w":��
��ଏ�
4����5�����b�K�X~a6r���R?s0ߞ�}���w�]^��%(��4�=^V�������襴�ȅO�CgP �����1�7s%(�7�9f�K��w6����o�_CQ����x�{L8����Z:��bĵ\H�'(g��j�[I%ג0�#,�AձQ�\n���@I�rx�}��@��n�*O� �׎k���nv��SH@���=
)�ճ�\�8�Y9��v \u��d�Nh{D�Ŀ+^��RZ�"6��1��������,��E�e��F���2w�ǵ%���&\m�r{
7yCyM��r����w(��`�a�x�|�Z`��Y��5\HP�oq]�1M{̻3�c_زf�Z$��yi6 ��6��Ȍ[���,�mz�VzVtI��D�<��
ky�#�O��.0�GH�Kg������z�X�>�=��\:�e���B�L���s��)6?ԠGC�ܤi�k��i�2K��I)�����٥�-L8f�P�m�����"��H`\�BO�R�fQ��~c�(t,-��c�\��k������zO��]���:S�S�QgA��c�a3��R!���q��k�����s���-�T2����o�������4q�O�Kj�o���"�[��� �J]���,$m����y^��ގ�t�Q�/y	�W�e~]��v#��a��8���qNrk�ulf\a�\�6tf�^G���W��ߨ�믧�V������S>d-���oN�k���^��VG/�GϻK/_�Ƈe9���۷er�;�]0�L"I���F;��K������ �	�yQ����80�X!\�!^�*���������1b��7ţ�Kb�l��1���M�)W����df�+�{��#h�w,��4-�����������&���`o�X?ޯg�yy�V�%-���?��U���1(ݭF!/*++̉.�b̓�q����������1�Y}����iJ�ΦQր{τ�yi�ƍw;�
(�2	���9�K���Ս]�u���6��ݏF7�����z�$�b�LP�
�ebfЋi )����D�.�q��f*��X�Wi��	�;Om?�7B�{�l�k�k��'�6����3v"�#]M�$A!��������-uB=xD��r9����CN�m������<~�HfM����f2�t�r�s�+1w�r�JYc�[�Y��o�kqeo�.�H�6vvN�soMOT��Y|"��D��|MGG�����U�5N�nl��%V�!�+����?�)ZI&	&��!����������&wՃ���f�E��
�	�R��m�M.���/^K޵D�:x#���[q"O���S�K�b^i"*��r�21OI���!�v�k������N#8��ՃUK��9)�yo�e�Q~i��)PIr�Y*����^mS�l�I4�LZ���ۿWV�W!���NYë��3���U��Q��O65�����|�sL�
�}+%���y?��ʙռ�%61O�B���F}Eyt ��-��1��3�L�<��h��˕۫&�+v��O�����k��D�Z*j�x���JNQL�5��q@>Bd�VX�d��oL�.ʢn�D�8o�6^Qe�����_t{��v%t�=�3�B�TAh�YdjmOfM:���x�R0+�K	�:E���K����sV�:ˣ��ѵi!��j�sg%⁔��X@��GO�I+�qѱk��ٳ���F��g��b��w��(���au=���}�aB��ɧC���3�,,��t߿/^<L]��zX�Hh���(�D��3jm�_<څ����]�|���/Ӟ�s�¾�(�N��R��hI�/.�A������f�sT��1��E���������r:=�o2?��5tx;!؆�Ή�4�${�[h��붘	��޳�Z���u��"��C�JE3��G������8p�O0��w:>�]������12�S��-�fzW���Ϯ�R�J����c�D�����w�ql�i�X�E6�^6���z&8�H$ڴ��3����#��mZ���D�Ԟ����'�~s����]G��.-��!ԗ@�b�\����v��ZOsxɾ WԌ��:$�M��z��Ɣ�؄��NkP�^k����њ1�����GM���^"�~�J+�Ո��hhQ��^�=q�zޘ�3x��W�*�۹
�~�~y}:I�Q?��Ǐ]�aR��y;<$O��d�!���}����W6w���������E_e
�w&5-����8��qވ�}kt;��_,�l��W�:�{۠�F�"�L�A�b�5�2�Rge��t�7;.�t�ѩ�iu#��*�G�YVo�^�W8k����I����ᠤ�Z�}D�@�/nK6G˙��@~t����Z`
E���r8ٶ��M�ϟ�8uՖ�t��R�3���h#��f��gR��|'���M?���G��-�[��w�H�::���8{AN ��WQ��X���>6u�n�o�r��DE�œ����'��|���9g��K�����}b�L��F+�/F%Y�dRO���@�����f&�Fc��x�6<������V�O��^I�z�-P�ð/.��\�$�D�!`�1w��|���"&9C;�
q4t��zs��b�hyӥ�����Vzn��½V��D��D\i%�(�%ֆtT�O�^�>DK&�s���9jS�0�I��8mCoSsH���|<&�|6*��Cq�Ԛ�!`�=??�w��Z8�e���J��6ssK�"��,�������v�>`��UP�]1��`g�Y�!�i���1Ȧ"���Hr��p�If�� ��M.���	>���8��B����;e:A��4��F&0[Ô�fX�F��x���H��U��T4�&T�_R�&�*1a�\)��D�[��r!x�ț����w37�k,����&ͭ�x�+KM�̺?R�\�f؉#^�ӱ\����_��~�S D�����o�I�QvZ@�[�K/���3���V���u���5G(5�`�����ܛ�[�<����&�]k������,@⋓�Z�v��gV�!����%Gm�Ɓ�mo���ƈ6����P�2��͟"�DU��V���#(�XXt��͕��$3�D�xNR1����g 5.�R�@�M��{Jcǃ���p6z&�vn	�;�۽T���1�
^u�-.�ҥa��r�I����Z:>Y����	�X~�m�s�uæD��͑m�p��\B  �ڛ��ԭ�Ol,��8���H�w"�|����ٹ[�f�3���R���:B�&e�n$ʗ��[(��Z;R�xj$@H!�"�pEz�9��yL�|��=���l�����CV���s�%x�sc``��,��/c�-�Y�BfM�2>i�C9���@xT]�`�����h�w=�[�1�b�J�G��'�ex��]�jH�i6��b8H-5��gk�>��_�Bo���k܄Ά�￭�*� ��R5�e*�
���b����,�'��[�I(�Dd���4��@��!87��ȫ�mL����p��fֈ��>��\�����ӸC�p0pPCQM$w��x�s������]�7��q�ղ��u�<��Y�No0	¯�	�|�0�����C�AﮘеKV�yi%�-F�U�0�l.����ϣ��.ٕN�B+���ڵ�|{;���	�>mʭ<���C}^�1X��P�2�|~#z���M�~FXK����aָ�K�gd.r�v�XU�n�yZ��5�������M'7��j%��$�/$**�5<2�	Q@	F�Q���c"�,������Cb�D^��-���(uA@i��b�|�B��i�;��b6G�[���W������a��4Q�������Q=�i�.c�����y���Yy�%=J5`���|C w�Ko������f�?�X�K�^e�d|a���~��J|fP���&�H4�ӣK������FLL�SSF��Ġ<�D�,O�4�C�g�i�W^�a6�U����W �|qĆ�HƗ0t�9�c����8����	V�覞^L��gu�f))+״}ګ���óP7�������&�\H�A �*:�h�� ݴ��c�|rܩ�Td#�����������&�pn��m�h]��3d��w��#�'v�.]���m�' ����I�l�Ye��f7��ɿ�t�[���q��f��B���k=���N"	OBx� �j��ı�)��~:^���T�~�sot��_�_��Q7Z{�~a�2j�dS��H�ia�^�?^������7w�&�Z��Y�(�8;;|�mZ���R#�z@m����ټ1��^������H���5������>�x�{�@��)f�������g��g&���aP�б�n��Xg�*��)���$�h$�eu�#�ѳe�qY#n�`g-l��n�M�G���>�K��p2/�'"���t�rrs��*�i�B٘�����O���[�����X(���Yp|�O2��Z�t��*2Q�[e��Z���~���S6�''����Ko�?���;��\>�I�Rb\����lK9�`q�M�G�`��*��T��-��z��.@��
:'c�k�#�o�F���~��'&\����S��` ���jEDc�Qmsd�d��sΟM�q��@@⦡}h2<���'qyόF�����N��?��W���lA�&�N�U�m[�9r�B��&S�}�ڼ�E	��;��3b��=4�E"�0�������T,�F���8�O{�Ւ-))�gt�<��;!��>C,���Ɖ�|"�/y��$|�svi�g��Mh�}���9I��{��)uyĀ���x�d4�x;"~�������^0�#�G�	K:�bk'+2~�+B��m�F�`���$�-X%�O|�` �Zʅu/��W�%Eu`z��C~Фd��aI(��(�L?���I���Ӟ��ea��y�������D<Fk��It��M�&�T�t8 ����,k��~�n3#�;G�)��`�Wn�4s���Ԋb���iD���������}� ݖ�����'��������OBK�=�D4>~4*�����Ћ��!�)D�ok�xHQ�2a��L_e2㞟�9�J��<�{���[��u�g?$��!s�q�z�|01�v��O`�y�/�@~�.0�8����?�P�Y��1@��8��C��g��W4�gMQ����u%�L!�-]=R�0p�O\:e>N�V����Mk�d2P;"��o�ˀ�˱tx��4�Xk���,�����**���������wa�z�iiּYKN���"^H�X�$$�P��׼|�}6�W7�`�!�qS!����\	��/�<���?�����8˾����<N�`�J�^o�H��r�t�^>����ȱK�惇@d&�v��R�3At1;�t@<n���/����ќ�[%�@P6����F�-iY�hӊ���w�yG�9���B}<R 8���}@�Z��#8����?���˷��(��聚x���dp�l�i?P�'<k1��ِ���AQg�P`�z��0�"8�w��p�8�=l�{�����u}�
�p��a�I"ִ�3�B+�d(���njK�d&�J`Աү�uڂ����?\��o޸Gf9���sY��u)k�1�>'sK��LF��a&��,��&6�Գ��&�w�Q�M`����%^'&Y&�{X����{0⨫�B�8$�V7�1����!����/��w�!Jք�|Muu�Lfۀ�z���ȥ����PZ}6���GX�O��i[�}��9�U���ճ̊�������}So߶9�A�+6g�����.�_0���4 �%�L�d������cK^�!��)�^13��LgӸ�ó>�`��V��ϚX����;��	�^9���CI#��`G�c�u�.g��DA_%��J�OZ`�K������Y{�'u��D�&��k)��ʇ��bA�"���j�x�^��|#o69�EEԐ�'i��<��C*�������451'u-�^|���^b�؞����_�
�}H��z�2�R��R�W����H��h�ѳ���`�ĭ7��.�r�����&���(��Q ������u2��nLǸ{݄�L��������=���4����"i�k���\�D��K�O�n4��&����ڌ���dO8�N�
nٯ�	ma�S�i�]��BHF���i�,?����L������x ޞ"��Pz�x7�BW\�A�$����23+ 9�]C1�Nn![�.aC�@m0a
��o�L[���3��/��q���0�K���@˱ܭ�U�x�D�
��߻)C_p��!��'u/�|U�DG���+��~I�&�'�U��>��1s	�|:�tSM��!Pv�AG����Q�Xė��Z�~��ޣ��E���:�>p����#N�	�w��ݣ�ʍ�-��*�:��Z��")�[�ʋ��;_A�ᇧc���+B�t���!oV����z��L�X��ւ�)�x��j�T:"��e���3J�Kl��`bQvR]�m�,2�:P=Ҍ�g��a�͑��W��ʵh�,u~|�7u>(T�)�yx����b=�p�~ʊ��.J����_S?���g2 �6�c���!]�c8Un�h�v�����^/�����ƘUL�r�M1�?�=�?��a2Ť�¸�}�W�5[��1���Z/�ߨ��⺆��T)l���}�,.���\{����P�3���gH�y�{}j��'c�&>q\�H��zs#ԥ��� D҂��]q/���ih�f�Y]]��s�ʕ,�L��sYl�����/B�啁!��"����<s��|b1�m_!��"�]/*�t]�?#�x������TT�5���w�]�T�y��=�}@�������yǙ[�����=�T�lRRR�����]`޳Ę�B�G�Ҍƞo,�_{���z<@K!f>��F�Ǣ��v�W�0R��D��)�[%���||P�2�W��"�=��n�r�fz+�ym����Ue�z����_��A�{rC��w����x�tA��&Z۬h4A&�N�s���[��|\I�ОA�a�ԘQ!:H*�$=r�ߝY��e���[̧��e�,BJ]]����Ȍj��^]�T�o�o)�zｳ��\�B�͗N�l�b������=�Ls��n8��5`�K�U8���ĩmn��Z�����:u܏w/=�V���X���+�Sg�w���?�t��H��|h���ǉ|'N��8�m�*�S��� �ێg��S�W�Z[��i��|����C��]ܟ�>�� �I��Q%�@t���ŭ��4�M������4��q�Wf���3t�zIZ���Q�\��
�ќ�[�Q��O�۳�"��bUЎe@H�Y������}��IO��K���ɡ����H�����T�BT6%K�����Mb����=f�B]�i�ה�D��aa���&ص�CN���e����6�L�~�k\��X�8y�+$�����qG��~%��[����؀yq".\ޛ�|d퉅io�
�jP9@k
M/ 6Ӆͅt>���1a�zPPQ�B�����l��;.Fx9COì���	3]�T_)�Ӌ)�g�P#
P-ߒd�`&���Q�0d�,2��J9�J�c�o�U�9T5�v��[�Ui?��đ��*S���(_����uz�L�k�8�8��}���o�^��տ*���~a�ʇg�t~�f���,'�-A��C�H\E²|��y�Q0U���D�?�?.𨗚����6�^�2�hS��:\�w��$���7���b� 5RT�� G��22������%=�|rI��D���$�x~��_X�ؓC9������w��<i�P�Z���'==�db	�<��}.�t����:��t���X;!vu㋑�K/��C���Yp+s�B(�F/�pT�S�����%^�V�o������D�|��e;s]xa�|��4�5����F���M1�u�'�ʹTa�~�{�I9u�04��%��
��M���
ŢaMLW3��UP�h��A�DSF���['w��k��P@k2����g�7Qb�m���{%Y�"%p��%��CL+ZK&��;Q��U,�i�ND���3��#�IiJ��8�{nN䝍��L/�ڷ�ۣ@%����7�O723U�m��hТ~-����岅���-G���ZL���t�t鹹��Ս����:1�0���o�3���̏yY�B��o��<=3$�9���pG�kT��2Q�ʓ ����d�V��@D�ܳ����՘�:'��ϥU�$�j��������J��*�=���W������q��-����y)y�h^.G(��K�ʖA�T����g欙�wŕ�U	���H0	]w�4��9�n>8IQ=�������kO��v��u���>&��^]S��U�;=�$�_�2(ͰeT�\J��*{4m��+�S�8��x��1d�w{����+�h�����m�Zƞ�V��ئ���qFR1�ѻ
��oQ`}圊�6_��j��e����@y��v�3RO��	Ϙ���f['��o��*�e��K��.P�1S�7��&�A�M����BMl'@A|JW�.b�rǇA�Ǧgr��٭Ǟ|�rèL4ֹ5mmp�0s�'0C_W�ۦ�Q	�i�ܤ�e�_�Ӡ7ک���2��vѱU��Sg��ك4&�� ���r2d�B\!�uuK��'�[�|E��.�)r��B�	to�G�U�z��?�=G���v	�&P f�S��2;}�� �Z\������A:F4��R�`��P��:��ԑp��	g4���'î�iZn���I�k���J�ŅD
��E:��x�Z "Q��;a��@�=4���kZgL�
@pmF�R�6�؏�+�~ᜍ��Q�Is�l��6DR����8�#�r��q�ub�ƹ�q������|�{������=9\��:�%�T��;k��ʳ*� �K��8��x�w������-�E������Gߘ�+��R�T�s����g�CAU�{Pd
������B�M�,9�ט�o���?
��D1i[�r�!��u�\�5,�����b�~:��ki�3��v�b�X�.R�����uW[��7���U�V�Q�Z�hfzj�ȁ,շ ��k�ڗ��C^�٘Ւf���T�ѿk�s�OK�\f�"]b�u>����{��T�BKw,�j���2k�_�M�PW����G��)Hz��n�M3���܇�7,V��K:��/+*u�TO�n]ua�6�C������nuM"�;�ys�x���L��PFǤ�@��*R� ��q��ZUKY�R��j~�x�f�4��XӪ�/yJLU޲5?C�S"�`�*�BS֩���_Ԡ��;q+tĴ�Z����*uT��F-��~�P�RZ��S}�Z�%������@����;9�]v�
��]���L�\u B�9�}g�\B���*�#���H^�Bb,x����%"������	�L���m��shi�i�I��o�]�q񃮬Z���m��+���e�_ۄ�?�?�#K���M(�S����Y�0�� �@MJB�B�������>�M�0���<;�o�wLN%OiG��Pט��.۵*�@���;�R�5�P�'������h� �P:)HU�N«�o�F)�y8ke _�m��qB� ��~yyEZ���k9Կ76sݵ�.��Tx���B��#���'9��P�v����qt6y\�f���{S���a�F>���?_����/�:��>��bt�N+���b������
@Be @��Z�8Ȼ���C\�d�)��M�=%m���<d=�un.�Qn�Q����h��c��2U����q�:���f����u"׼�Z��<�|K|}��"���oڱz��
5��͒�\�a��~��bq�K/A�����\�r"���;�S�(�\���6��ނ_-8��WD�ɭݨ0�hgT��͹�����0�x��<��R<u��m��O۴@�_솢��r��	��͘�O�^���*L�?���.��f&��u"�vh�h�dM3��w��{�CFc����H����>:2��U	����c��.d,�-`�[��1��DJ�Ө��D[���IA� q40�M��z��|"E:��i���7��ë�!K>�X�6�����/K��c?�$Z�d����vm�=�^pnQ�|A`�%�Q+�Z�&����U��]1r�2j�/^(�s�Xޞy�+�;p�V�����>A�S8=u����߭+MYU�<ۥ� 	��+���,�[�I��'�t�K��u]��v��U�����w��m�ݵ~~?���u�4b)���o�Cz��QjPGu�dԤ��ցn�y��i�w�15�Ly���T�t�:�q�s���Z�y��k6���f��A�Pw�>���2���)�3�E�elꨁ���6�u_eQ4����|�j�U'��Cbb���F���Zqu�	Br&H�&
@��F��+��+��+ެz=���E����D���~�}%�u���U�y��͋%�2ͬ���C�!6�B?XW�и�ԭbx��`�u���J(��)i��A�K�$������5"e��I�/n���z��+���c�de`e�J���o����l��HcT~����o�Qn{� 5c�9��E(���1o�S_�\Р!��1S}�qǷ�wх7��r]6I�_ބT]����WXo�NO���:a�MHBr�f���Os�H'�);�ȍ�5ǁ�!��̝w�/��/8fֻ;�N��6��s7���hBǧ��*��8��i��Ӆ5?Kj|�{����!M ��S��������E�� ���7��>�R�K^�A:�u��-�'8{� �;ߚ԰󌹖�u)}�~uMQ+�z8U޻cO�[�t���K2M������R��v����G��I"��)[��Q�LB^->4מ�i`R�T��qչ�ݳ9����BH��GY��)}���/�����5���,��!����� Y��(k2�����'?�ꭔ��n�۲E*]�WS��մ����?ۮi�@�����/���sz��(,k��(m@+e"-�*	@P�-gVTJ0M�%E��Ad���#�@�,�cϒ��6�ݔ����AG�`��zx��u�~�xW���߆q&"^�.v�C�b\�Ϳ-��?���Sʴ�6) ���T�,�U�
��V(�W2�#-UOo��'ԓ�*�#�h�\0�-q%wk�H�_���Wld����bJ~������7�h� $MF|��usk�׋튏���e*�{u���b��~��;����0C]I�x�T5�7�ꓨ*���)r(�#c�xZ�1�f<㏨Z��g���`��?B0��Q����H��c��.bM�L
F< q��>k%����^�"����n.���#�k�BS�2&�5ʭ�4�x����M�,����j�VL���NTMil����;������{�nL��	��7q�?��H���?�7̶d�����%1��y��cט�G���q	�R��ϼ�A� �HF\�((�;+K��h�}��Y.�0y� ��c3�����rM8��'3%F��M���e��i�^6T�Z�u�h�x�3ʹ%z�3鉟���v�޽�ȟkr�+��|}=�@(U�S��Ko�/b���u��`s���T�����|�v���{ t�k�X�.9^bY�ĠF�,���w�I@�C�a|�E��s����D���	�np�:|{�KLYu�ib-d}x�d�F�C�������۬/��|��a�)#$˹��L3V���׭���J��u��4��&����)��n���	+�;`5�2�uc�Io[_���p��&�*Wv!:o�c�n�i��hR�~��K� ����f:E�vT�}�4��a��I�}������#�8��m�=.�R��h��0+��N�%�ښdv�a�����F5�E$�-�	B8��D���S/�@	H�@��Q���:�x��$��E�g``��Ƶ�(yjnџ:O[��?��k��	]�����vA��eE�2LG|,����חA�CG1�m��*Y��5�cX�jS������>��I`�����p_�˕�O�	onb�`EE����3�i�{�wn�Zy� ϛ��1\�\�����M2�{u��A.ˤB���>B�����tz��Ͻ_�����`9��wtLl����x�Wq�0�-g|�Ğ�I�w��[f�ۣY-w���*��q�A0��&��y�l٢���.i��"5�u-�x"��	b̌��@`c��۵DA�����m��}�R�g��JZ��}�#<�8�D�ڏ���w�����G�+Ւ���6Ȇ��M�$�#L���|ɡ*-��(�*o����ˋQ(1{_���=ȝ�Gvμ�e�pJ��kC-�o��J� q�=���USG�hA55���j��cN�(�g����-K���j�y{}��g�}�b�]tץh�B�^��qF8�A/&!W��T��>�K�N�k��� �v����mS]}��)���YTΉ�9Jsߤ�\� ��8�`h"ӎ���}��|Ӳ�΁�6������B��펉2�x��s�
����\c��"�W�y��e����2�:/������8�R���D���H��4VR8�ˑ�E˖f�g�M����A>�x'������'�������_��{zz���@���|�i��"<��P7�b�7S}�Sx|{��
�,ЃN�4b��t��u�����k�8�U�W8�q9x/.�	k����j5)�M�>mWu��9�C�_�x�j�B�Ad<ޞ��0e�E��7f��Ѣ�|FN�dolmR:ǘ}�,��ὔ��u:��u����,Z���ȵ�nά���w�9%s�	a^QW":�H=o��0�W�b5�|��'fT@ͺ^�a_yu{���6su[�RY���8�18�$���E ���Ҡ�ǭ?��˵@J������z#�H����y�b��ԚŪ̔�]�M�Y� djmM�j[�*VE�NU�$�����s�M;ɀ���e����%��4�9�����2Qqy�4�h՟�ɔO�Bg������NA4a�F�`</'�v�$��B%Z���<��|�y�h���8�|bv>��\�+�CP�w�b��,�9L�M�i�d��T�W�!���B[��z yS���>tygW��-�W�a�k���_r�:��6�����T�R�4���JtRtI����`o�u�g l��g��g�{����x�Xz�_Ww�B����2b�NEK*T�3�W�)O9Q�8W$�ۅ�wsC?��#Ӳa�Txl��YOG����~��އx���/��8�a�����<ދ���L�r����oWNsr��;�<���Z|5o+�
��z��P'�_�~	��1�IE,�G����j
$�\��dT[p4��=#�q�;��ĆƓ���]�Վ�W�1�,�RR�Z�d�7��р��{�.D���~�"%���!��@�ޚ,��Jя�L
ԙ�x�5�l"�A�O��0��_3)��>F���y��o[DZ]�0�;K��R1F��r�t~��@�0�RHQM�JSCu?s�3y� �
����QB	2FP��u>���Ğ�9�v�o9�e#a�8���e[iOʈT/�gTҔ�����o͍�W�G�@HD#[�C�;��*��.���H�ib�w�L�rL o~�5�/��[��ܔ*x&� �v�����"��_b����)���+��o\����[�m7�ܦ��w=������h�=�軼�@��\��vα��q�];���g�Z���6u�q�ݡ.[� �i��㻿U�y�zI+��T������h�7. L4V
�̌�Q�|���#�q��}����ƃ%αT(բ�l�[N<+W�:-n�[�����Ao��f�ĺ?��H�a��O2R'�շR*+�6�@�#���SS#^q���	a�� �M������g�Jtu�����h�;x�R�P�@P��{��y�uO��8EȖ���:?M^����S����%���_�Р�ә��H����8Lȶ�J^ �:J7R��z<JjZs#ɲ���m�.�$�~��l�nM��m���S;?���<6�Iܵ9��}����Dħ���8���*��~!����ٝӿ�USQ��ǳ�}�)�%����+�������}���H��·�'�
�u�W�'/KJK<"��^�Q2���R�gd�k2r���A��С}�\6�J�4�� ���K�x�|#�I�y2��7Cf:�7론���+��W��rc���W5�{GWP�M���]�˞�wRv�o�֑��`.O���Vy������r!b{���[�Ӈ�Ӈ��;F��=L���6@��g��bH�i�<i��^��¤]0�Ă������\��kjj��εB��^ #>��#j�����r�Qs0�~װJ�WROB"T��`�_>E�yy�����gP$ҭ��Y�6�r�ـD֧�=槓&Ѯt��W����򁇀�9G��Z���8�[*���� :&5���Z���\���s�! �����?��hh����z�V|Y^��[2�4_�^��*P@������w��N���4Y��(��K$�'�U����CO�*��=U��)�,mf���c+�����O�≍�X��)�яC���=>[���Ҏ5K{�^���fR6k5Mҽ�sF��e;zq���h�l~	|�O-�$cݫ�>\��_��m�^G�z�J#C#�iJ>r$ǩeꠖ���Y{v�Y�PgP�F�B�E��"a+��>wi���;�l�La� Qը^eӆ��H����|3,�eB��>~�RjA�>:���o����w CF�pLx�W�IUiu<��z�a?�~�z\J^r嬑�sw�|ʲ�����מZ��`�=�3n�}"��ū^��V�^Zgo���n�53�z�dY�)d��?��b1a�q��$m��멆
ט���ӱ�koּg�=\ ڧJl��qȶ���x�Dĭ�Ϧ�'��hq9��@zx/��e
�5	@�/`�Os�0�m���7����%�����H���r�U�m�-U��=˕V0��s�(߃H
#�'s��=zgg|*J̔��8{�4��f=��|j����Uͤ���`]/��r�
ʒ��S��Aj掯�J��Y�:��z����dˌ%�C���7O��9Q^)q�?J:�@���p�fiG67Gx��Z$��y?0�yo�f� �)#�7�"55R��G��ԄC!`%=�?TG�'�4��` 2j��`�ݺ��ں�(x����uz
ɮ��>�Q_<���Ĭ=�XL����M�F-�K�6	����i���]Mk�,yC|"!��<�����v�|�8��z�*���9��e�~�sO���T}���GĘ�7���ל��~Ep�9�B[⁭g�]��&��۞����	�wc��c�c�׭�Ԍ
�=J�4�<���ud��­���]��o:�~#�1���?�｟@~�/�pi���G�����H�<��H�;��z��|�2�8��0˲J�E)��*��� �/M^�P���=?Ɖ��8o43���﹞�	�|�%����i�m�����,�Hm�j$M�֥S�Gn �zMH������V��cd��<��Pu�0O�c��s�}>�����pH�38j
�є*x������衈���s�A�h4�T$N2_�.�����,0R}�t����);h�bp{��r��V]��D�7��&�J���u87�?q���ScH��L�K�@���c[�I 	p�&+�k��T��A,Ő�9�<���L[�4�Ζ;Ef���=O�@�*);u��o�?�ؿ>.q',��'0�W��c-��m���J��̮EQ�= �E(���M���I��ы?Ǿ����k��lq�G���p2�nԿa����$j��Dh������1q�����h#��Nz/�����p��{��"�
K/�t�4Hw,K#²4H��t�t7H7�tw��tKww׻~����̝�<�s�{g&��`��e M�>ڍ���Y������=�{�||�xu��[���ԕd׸B�4�2���0P°�,K	n	R�'#�8(����Cbe�R��;O]JmebY��m��٭`����~%�	�F�A��#�Z���ZC*�'4�%��w��JL��w��壪�a�Sw��!���:��r�|~�"�$�#��H�'2��u�����p������a��SR���G���<�@ߨe٦�s8���Ҡ��=jd��u�d�f��׈��-Ut�˧�ү���D�f�M��iM��?����G����2-������r��; FB�Y�o���k�XF�V����͈�>��5�?��g����qX6&W��,��c�N�0���t?�|z�8�O����:�*�2 �s�`<��zd^��2�A���� ��l��"�R%x9��~�C 1��ֳ���\�.攻UN~;T��}㜯��΅��J�������x'%***3K���i��/�?�5��o�Mϩ��oF���V?7�dy����Yz��}#��Q-�D|������}	�jq�TêWrj�Yk��o���R�|�,���d�1�7۶��m>Q��}t;���l.��%����}L��� ��l�S{��qd���!��l���vok��iG��?@�Ǌ?U�#��}�n�Wi���ME<�9�mTon	N��/�N�䎖3F��G*����F�wy�.�*����r���+�W{g��y����8ڧ�&�����J��G�Z�G�)��L_|��E���H��?��� ����������;L��u����ߪ
�}��m~�n��s&k�4a�[Pݢ'Y�(ԃY؄;K��aY1ʹ���}�D.�]��+�]�X�h��q�@.!"k��w���A��*Ӷ�^�`o�C�Z���P���?G%Z߉�d�}M��&�g�2�@xHh�|�p^�YV�*E^ &
���J�9��W]-�!�As�WHaÿ��1V-��i!��fN�=$s�r�d��͝�F}�$//�&,1��+{�IF�ҍ�tN�ov��C1^>����OY�b�WZ6~�=����=�kb���Pcq*׳v
��K'��������깮��l���j�+q�ʀ��J.F��U��⬨S(���b��� �� ���?��=|N]F�:G��E��J�AZA�{�^0��j�Ām�u1	��R���d�̜��k������h~L+�^� tT��\�����Im�M;�W�*�\�#������Y�)Yr$�}���2֫{�S&l��6K�>���M����&G�Ls���4Ϳ�6�w�C��4W���FҮ���؛�)Ed)	�JT��؇e�F\���t%s�j!.R��[�����y�i��K�-��ٷ�j�-�ĉ:�������n%w�0[qLb�;�kT*��h�\,���|�u�.!���P{�����]D��2�F�E����u7N�]��>5�8�6��)C;;����o8���nowQ���]2����j�s���n�p)��!���:��9��\0S�-�(*C4�˗�������G�O# �+��箇���$�#Ϩ�[$�<FQ$����\�^��B3It����cpK�	�z6��^�B�j�Er�e8�)YS�a�b���vĚ\;a
]���ՀD_y���$Bu�ALV��1�m����$ T�B6����W�
P4:;9 %ڼw~Ĥ�z^7�13~���'Xk��tȔ�٧V�%��;7�rgӋ[*g�:9ၥr��L�V�i��g�Q���}���`����^0�DL"1�T�� �r��l�4������h-7��.&�Sy�18����ZQ�2XVr�ɪĭ%.ssb>B��]�F�=��y�����O�qo������g�`t:���|d�A�F��}��D(Z��y�P�`OuO�Ք
u¤=5j�Z;��K9TNqR��I�#���H���r�tdT	�l!�ᐭ�~�\5n�j�A*iR)P-�u�񧀣P��h��(X,K��W��2<��pi���[��݁d03^((	V����K$7^!�l*�����!I<S�������m�Թb?l��e���;������3y�[�8�<�j,y3���Uu��h��D7�w�H�jA0����QX�����b�W1Z#CY	�|�^(��+ji?��I�0]?O�5�~9*}�ZcRb�w&���&�Q6,�;Wap��s� ���|�&:A�֥[50L�Ұ紇��c�D�f~����-�����h��(���Z!�v�a�y_��o�f�(M1�CX)K���a3(�H3���ZiN�gP�X���+��9�9���)uxF3B�ؼGQ��q��eXR��Y���D��3�TKd�ֵ����k;���g����P_� �vc+w�
X9�N��#*����Q#�a^�"\�����8:^˙iEE���n��3?�o�3��ǟ�Uک�N	��
�-��E��Iҋ��t��&�$��̧��"��qAA�؍B�2��WקG�:
��#�fe&�Uo������&�q������A�<�K�I�]�qp]���`��-�#k�kV�
E�-�*�{��|OECg#�%�C�¦̥�G�#�7��бF�Y|�Y*�{� �����ܼ�7r��wv90;sX3)�&��}9����u��ԢR0�K�G�A�S�]��X�N�����<(�����������m��G����{��'�sk�*�`��{">�p��<�����l���Գ�4�Ⳗ��FD}d�?�[}G<�`��+��WMSv�늺�������C����Z�r�A�n�Խ���bhB�Ş$n��Z�=	����~�i>�o�p�\�͉�K��M��#�Z�u�݁_uAGך%3'���(��E��՗W����;|m'D�C4TZK����~��Ƭ�G���C�8��{��N�2`%���~��Ǚ� #��_�i��zޟT��ۿZ�;�U��e���=�^�"�DOO�p}��.���@�C>D��f�S��ʧ��r�~,���}�ׯ�3z^�>w8n��Թ~Y��5��ϱ�}��|1$�p��?�x�@��F�e=�K��\54�u�P�����"/����Ul�C�M(4㢸��s�+?�y+"-�sL���֮�,%�ӣ�M����>o�����N*;�U�)H|� �}��~��Կ9uY�2��/y��Ji^��<�٩ذo��2m���FO��=����I�s[
��b>m�����ܶf�:Z���9ST��bnbQ}������N^�0N�B(0��8��hӽ.��ݟ���P<VZ�7�%�⬅ژ�-C�g>�L�?����:Zu��$<�lV�Fzwx;��a ��d���y��\Lp��P�կT�殮��a���Z�>"bܜ'
V1o�o�8o5_��cz@;�@�z<aS��E�ņ=_�����/_��Mo!��ߩ;��1��i%T�UKs��t;�?�*P3��xX��NV��V�1��&7�!:�BC"σ�__�NFK�]�ɔCb�Aq��a^V	~��8�*v���9��eҶ��#�{�WQ>oeY[��K��H�M��%�q8Eڶ�zg���w~*���Gd����w,�v�`�B�<�b.3��M6Bɫo���9�t!7���2�۞�E]mp:����H.vT~ƣ�	㌜�\��!��A0�-\BB����c��b�Z�j���LD��y2�<� �&����9���R*�f�x�z�P(E�a��E�ٲ���w`��;ۍG2V�Tg��о�U_����凭�=��5޹�7�j��4��cozߓM/�c�u��b�����S����,��`ڰ%d�^��ƷIr�
��HU�"l��V�0�Zᘠ��#�/W{�:&20Z�[а�Z�[u1��܊�rf���"E�m�������'����?�\Ѻ�!�ȸ��"�y�(.��V����/���Du���w����/��A2򴱷����O6V��~�מp8422� e�;�on#��l=.sǘ��J˓E�nV�O�rj���}���Ir�=�ۍ޶{w�玴I����O���1����r��j��x���H�R���b�A���<�K>�
?�g��4
-��Q�)����wP�#i�ƺ����ZDq���.�����PT.m��7�]�+.��]��r�-+�%O� �R�,���v���R��,a�euϲts���4k��lg=2�w �2,����l�������Pcd' eQ��A�_��[;�X����D��ߌǡ�%��QO�gt�NYX:�eq]�r�Yy�'[ݲ]�ks(|�`�Xr&�H.���NT���qI
	��Ȣ�rC�,�$��+��Z2�/�n`�&:�J�\��Y|�4�����t���U�EN'/e�BE7��"�՗�Pf��@AX_17ze4�D�~m�:�>�x���4�^>���Mn���؏�°�0��h�8`����Ô��â=�������C$���� ������[�ς��䌅lW��q1���s��(�s)�IGV��+T��6n'���-*`e�d	6�v5ҥl�������oSC���uӪ$��.��~��S����_,�ψm�ۗ�D�]X}S�֛31�/����c].B��%�wm��a�AH��aXe$�kO�g�/�O1 �Kƴ�]��מ��O���(E��/��TO���T�1]^"r^j�̸���ݯ$��������������bI"K�`���n�T�S�v&k�o�S�fu��;/��mA����gAL�����җ,3fZv0�d��i����Ç�#�U����5�� �-,w"�c�\8�ʓ! V&%{ꗹ]����ٮ�v���vn8e�[�_C����UӟY���s|"f�3]F���c�<�L�W�g�@��W��)Ԡ��!�_ax�\�x7�J^��ͷ�&��f8M�N�v�=Q�L����c��S1�����*����r_���* B���P��얲��n�%���1�����p`a	�����Ш�Y"5��*�o䙋G�3{�JJT~��l���-��S˞x,+d�o��#�å��2S�d�{ٞ�h�Et��r�ɫ!,Vߚ^�n1�MRH�g4mǩ��ޏ2�0��竲�i�֑��aɊ,��m#A$�ϴ��8"&4q��jsv������lc�:NNw	Q_��7������3T�? 6N���a��HFCpo�d���Qse7,ζ�S�PVJu���v`� �⃔�� 9p�{l+9:O0��G��N�q���6�'��U���F��{U�YQ�kB ��b5��<�v�m�����פ9B?P��a,D)#���4���_C&Q������R��_�_��n���Gp!yH��t&��jm�CJz�=^�=0���t�s�=Ϥܤ����'�0�� �m��6�G�(��<J�7�hy�V��h6}GK$H�A5����f�Y�����~T:��e��:�4�Ncf9{���;�L�R�UO��.K�QhR�����0e	�8AQ��Z�i�{1�E����<�M���� ��#��A��Y�(���7���c��B��9J�C��q�x�C��Y�7+�����Dl��`�R�		&����#�DZ�J��%�;k��տ*ǰ)d��$[
wkn�Jَ�/��ì�
o��d2�?��KOJ�`.���l����]���p�4�5ml��u�פ��u�'Iz�HNV�*����ֹ}��ӑS<�n^.�:�;%O
p',I���d����p��
V����&Py�(@���j���HX�j!CV�X8����u4��N���Zsϧ4���r��"r>B�)�0?�?�,���[��!3��
����F��b��qa_�5��,='�P6���j`Ɔ�p��;;��2˓j���N
�`f'zR�j����:�c��sL�8���C������~�>r��kI�X06� ��~�\7̽���[�@�GʖI�ُ�dv7a|�_�g޶X���n͵���wQ��s��J���2��}�VI�FŠ�����V`/��	�L�p��Z��7�]��W�O��Kd������!������~^U�fA�𬹾�J�沗�P1ũ <��m󴳔�S'�T��P��eD��Nt���Q��<)�$0�Y�K��J<B��7$ "(���C�Ho빯�C�`4�y�%p���vɄd�$u���Ur�ٺ��G��ܔ��(e�Q�H�&��n ��&6Dz����M'0��ח:5_����]3�gҞ���Z&A��E��ys��d��_�.�����Pe�4�?i}A�]��	�aߧ(�v�Rh��M��M8��ϙ��<!˓���8W�l�������]���8�D++ū����'@��� B�[��]�ý�q��?zQ��3�fC�)*��D��3T킓���Ǉ��g�a�ׅ���WY��ڰ5=����aXK��FA�����I��a:�!53A4���L4���x�+��n��g�R�A>ü�GDQ�ƪ�@��`#�����]E^��R[&)g���ݰ8Ø�.徲[I�S�DP�Z�_�4����1��mbߊ���z���PWi}�^z{�淈NK2���K�?i����t��ƦԶ f!V��C�D~�����=��� ���B*��n�;�B(_�M�9ž�#|�Դϥd	6��.Ɉ����6_p�=^~�:����}�*���yMfln�?0�X��e�%�a![�Gy8�\�U�shG�{4`)i��W���H;�|�rf_�8'w��TݢzҪ]4U����|b��t���F�������RM��o�P%��������)?�[��P�1��,S���~�j��{�u#?��7۵�;��ۃ+K���������ah�5��db�ݳ�T�X~���u�������{�8U�T����$A��ʗ�e�Iw�FobF���E�fJ`ME-{i�o�=(j�&ƀ뒷^k���f�b�v�y�O���o� �!x��Y�6��Z�Z2����G���h� 2WajI�&�Ն�fV���r8r�>;��N�7�W3���j�u�-��!�6(K?>2�?�����KJ�GM
ZXNd1���v�3`�%;E��.�vEC�]�L)o���5���0]9��5���Bs��Y����k����Ũ����|@M�4T*�ie��L���q���8��X�L����Gq0f3m~����^hHA�<i��yY����ik�M��gx,��a;T90�WV�R�`�`��`����V�$����PP��"��N
�&����M^�9�ߴ�\.�����wlL�}��ą���	�ܻ�ߴ�gbA�zϗ�D���i"A�T]3���۴���DGf0Ű��YB��
S<h�1qڡ�
��D�H��1=4>2��kN�r#�m���Sq{W���q��/�g����_{b��J֊��^1F�/�R��R����g���a���e0�K7747F�'~fu�o��@��Ò��ȹ�'������N��24�
�������8
G\u-��3�8��!��\)�P`��ƥ����������5}Ҭ�X߸i����?g�� t:�����& Z�뭰R݂��MD���Å�
�k��r�s���ѱ��w5�[��ٗo�S�)Qz`��Gcb�I��F���~���>Xb@���&i�&6�a�7y���cE�#����=6���������4g���=I�1&���O����U ��w����df���'QJ��7�!�����'�YF����F�����V�D�嬖jC}���C���N��wwK2�v�[X�wb8܌��"��w8/��~�z��|�x;�����#��8nQ�=#Ô� Ӗ>�.�H�y:�
�@�gn�5�ܷ=ߧ6�3KKC�'��4���oK����l<5��c�'�@�a��5W�;Q��ih���(�ś2ʯ��??!�ͮz�����?�z?`O	�WD����VC�;���~�.
8����M�|��ܾԝ���C���F��h�G�e�$��O�䠍f����`TȇJ'J�s��{?�-�o��:��yl��nY��+�cj�t�1�D!�qrV�I|j��h����&SD_���C��|~��`�]:/7X���E�ߞFY��f����ײπI��l�oC��!O���n�u�4�P�����7�3�>�o��ᶄ��'��i��ޗ�i�F4�+�����T�^V�`^���j�]�=00<�A���ՙ��N�!�VI��G9q�+��"����XYE�8�\������>����\Y-�[P�mG��D�c�����d��J�u�� 9����8%n(}���?�����=?���
_�a�Z��"=m�<�x^������Uo����3 猑�P��b��<mW? ���׷[-P�p�F��������ل�)2
��+��%��$��Y9sw�-|��Çv��,3Қ��nG<�CY��LĒ�Z�ol��3�����H��}����-͈�t%Fc��� Q�:Of����)�>^�h�lf�8о>�<�<��IhWmk���v��� u�ħcq�<�Oe���	oKLꕠor���a��tr��l�yx���~q.�Խ�R����UYQ��$���Q>����_�E��wB�[8O��O���1�5K޿�N@\ ��oL D<T����9��t S0�C�^���b�'*��|�t}����E����q	�߈ĹX_�'@Q2ޣr���}v�Qn@?pP�Hˎ�T`�K-r,wu�X~z��?����9��[��Z�����%��MMv�A�:!�4\��ABOJ�]xt���bP� 4�����<���½�*/*C�?
=��_����>�Qp^I]/���v*����c��Jz������E����zvЏ���-���������K���F��t�����f�$�@���A�Ĺ�%=�E�����տ<�릣���S�$��PC��,���,$�t�3U�x�����������ݵMWh�[���D���m�#��܄�����E2@�`0N��,�*�:��LT�H��}�e��q��l�eugP�>�>�g@����Cm�Z�1�:Y��j�[��Չ�����<j�,�����v�j�t����5r�{��x���\7a 77�(�7rJ\�B�y̟wxךt��.f5_|�ߛ�nkn�|z�q˥�Q ���g�Y��,vc#+'��n�\�ѱѡ71�m�;�8-�U%OD��Ld<H��O~�k}ŦJDb洝���_�;Ѭ���_nX4�5�{v`؂X�ˆ��(�����E�^P �b��i���䵤��)��J�=�FW���nK�����6�y��	����>��;/τ���Rs#����s���:G�b��
�FϋZ�ח�t�cGE�%��c�x� x.儲�Dȼ�&��y����������(a�#�#q��W�]E<j�g���2�J��3��Z���0���E��C�^)Ͼ�E|�2�יd�>�7e�ޞ���z;l�p�TV05���a��IGay�⣒ӱӮC� ��3OL�/! �='�bf��,�jp��wύEϤ�c�3=�!AޯY�(��
�ZZ-�����K`;�1�'���&*�$�WF��I�u��H]�05��`���x#�*?��3�Ozm����&FLL�ҏ�f��M�לRL�|�٠%6�np >҉�����&�J��3
������'9
j쒞s�_��$�BB
z���X?�P899���+��� ���!y�0�B4`��Li|M矇��W���?�i��K��a��|w�+���9Х屁$��%�h���*��?M�������Zz'Xl^륱7�?�GIY��[a-4
'r���u���d1�S NH�D�G⾞k��"<�[U�9v��9��
}�0,jq}��hҥ(�{D�5{�� ��H�L��NG��3�6��H�	7q[��".�c��Yr�f܆��r�����n'���S:��9W��\�����M�
)���-�A��G��J�ۉd����&�l��\���/���]�2�e8to�ꔎh����l��gJu93n�ӯ;�?�6^J��k<,�ܖ{dܚ$>���|��B���G$�(W���EdBRe�SK�j|
C���		�$�?��;kms�s��X�#��w8"F/
N��:4,
�
h�Oo�}
Qˣ�6<��&�$�yS��_>n�?U�7� �`SyD5�gGW��F�}�Q��֏:�� �����˅g*�t�AyZ�w���2����U4�t�%�n=���b��
�f���o�C��]�܍Q%f45�o)���@�e')#����eXϹ`��f@,���� V���E��/����ev�؛
L�%9�v2#���Y��^#�҆��*Q`��+�"Ĕ��U��-����jS�Jފ�f�<76r������d�XS�q�:�&zG֠^����6�w|ܛ\�O$�T#�BEP@)�B!{b��Ld��:��v�)�0�Y�=g�r�Rl��W���{��1ę�Ll�ܛn~��lV�O��R�,Vr�FU�dS'�R�íT�%���NS� �^�Ւ� 8Z�<�� �����v{~���� %���y����1��ճ�8]w����������}?���-T�����P1P����]o���W�C�h�0��s&!܎�!�Ao������2�-���2���:����4�]�����T]rRQ�;�ټ�1��pn��lv�d.�p�y9� vی�KY�X��Y�Z��ao��#t�ǥ-��g�����j���4�X�m����)�I�NǢ�^��ge%V���b����9�S!_7v�8M-	g.%��e�4T�3��<�bNhae�%L�q��l\C���$�𻮽��|���x�%Z����t
�n����P{��Vf	gDs."&���-@�\�;B�x����>�p�Bp�D��Ss3�Ͼ�PMKf��a����b�������sh�ӻ�������'�ֳ[LB1�ϸ��c�1�~���1���LQ� MH16��\�,7�;I�Ό餄] ��z��T~�|�VŐU��u��Pz�5��kݧ�������.�AU�ܴ�/�����+�)HA����P���/Pikȅ��Ѝ>�7�7�G�x���`��%Z��Z߹h�H��f��o��I���~h4x�Y��r/�oH�g��}���E��Y)бѯ��߯<ZB�V$W����p%���F�����a�q�����5V �'מ��S|^��9)�D093�����o��bͪ�I��>Z�eىҳ=��>�F�qQ�/�,�$��qM5 �(\��X��
�@��`��0Q��i�܀؈����{�j�����x"�F�]��!�o�C=���xXl��n�SGǀ�g��$*V�|U~P�P��ʄ�Ҍ\����&�'�J�̆�vAm�z&��~������I��!��^�U,��y2Ѭ�Q���0��F�(�0ׂuBBB�D\u��pk��w�7vU3σ����TE�)��Bjje��P1��	oK6�|�"�5;%�Z�>�L�z¥#To��x���N�?n�o���96�fhU&�]�Ӥ�p}�!�P��S�D7F�4��ȯ\<e>�h�LP]cftb�(���c%`�eq��B?�Z�}���~?�C��?��yWQgkT:&�暬�'�%�{�%di�<�I�*nQI�����G3����+���D������m4�Z{�v��M�?�*���������H4���%{pm[%��/S�H�%�����Y��w�aZڼ+��^X1��C�[��c���W���<�m&����,���M�O�ߍ��No�^6b>N���
�
�m�,�,�ܻ<�𷉓�J��?����I)2r���@tva����\�H�&��4@U�3�@8렦��������_P@H�v�jdk��5��7I���|/����~�^��>oRҒTy��	�5�ig?�R��6����U���%fk��[�^
&*�R ��Y���r��_a>t iCOt�#X���q~�)q�?x�l�n�?��`%��B6~׉�`mȌ`��$�4Ƴ�,uA']
`cS,���嶜>�,H��=,7�C�ɽ���Y�bm���a�."f�4�E�H���K�?���eDH`$��|O�=zr�*���a���h��h����%98ݎ"~���o=Ƒ�
�����V/oN^�����:(�B	t�Z>�� ���.�e��[4SLl��Y��"����yB���4Y���YoJ�^r��!k��[���Or_�4h�Om�)5�j�_Q#!���Jb�-�A�
U�&�er͌�.�ښ�ҫ�W���{W ���R(��я�U�5�t���%�Y���<�m�"):4�ܛ����D��)�~�>�^�(�\��Y���7�����Q�Zu�P���u���X%�0q'Ey̾7*uu=H�Z��
�TW\Ib$2~*��x����e�?f�����H��
NWi�_�O�qCT!a�~�,�ɪ� 22S��Q�D�tt�0X���Q(Tj����0��_�."9�Үޓ*�7'9?d��\�wv�?*���=Zz�/,Sut�~�E	>ag$����a�����[���T�a"a����
��c�/^��v���og_/ɴ��6�5��DQU�cn5j9�Zz�
i�^{�e,��MȽl�zq�IQ�f���־|.7*���U1�X2�G��h�r7�6�f���M�灦e)O���	�M�2QI�֨���Y>D����{NA�A��l�S��y��"���)������!j��B�$;ⲍ�+.7�֌<�xG�+�����<<"��z(<�He?�=�T�j�5��TJ��Z����lMlR!\�p�v���Q&��~�Ϭ�!��x��)�p�*��y�a���k]oO��$9�d��fKN�?MR�-i_�WD�"�Fi�u3�L��h�H�o8Ӥ�	�m��p�Ysw������^�	wD��X��W�j�62���U�e`�w��{�:w�*J��8��e8MU�YX\�x 8���w����N�͇<�P�(8֯�0m����4��(x+�t8�f���Cn8�MҘb��89I��F��!�=������(��sӋ%)ƥiJ�[�"�/�#��T8*���=�.B��AN3MAk/C�q����65?Ё��:����-��r�����kRƕ�=��!�H�h���0&~ON�.+��o=�Ou^�M�r&[-�S{8;������z����`���g;����M���pw^��R~��,���o�_[z��� ��=d���>��nN��)]��պ�dɱ8��gU",��=˷�y��Bz	��X�71lًG_��č��C$�ю�����i��5�����9��d�[qrut�1�X	~�T�5����ټ�%RMY3_�	E0򉈒�|�����F"�Y�E-�f��H7�F*��M��*����ړ�=�$���\S�������Cj`y����N&&&�NM�y��P({��xox<�>������{9��uPk�Ӯ����0M��j���hB�z�8I�j��B�rJX�5�&���2b��6�h���W��%������z�*i_yE,�G�و��*��^˻m�(`P�S���3I���Q]����|.��,Z�����H��ҍB��.��w%��;�L��#�,A�7�����Q ��JhZ�?���Ԉ��c	bi���^��X nА]v��B�}�f٭����)�7��t(��ݍmvu/�����d��)x�����҃`9]��Z2~�4[��^�I���u4G�z	����ȹ�3��������o��^����t��L����w��7�"-W��̎�!�����H������F[�= \�xЖ�;DK�O-���!`�������u�����@m��.;o�Cv�����T�ں�'bYq�jvT�� �8$��T�I�!�������G��QMGe3�4}��=�WG�u�F��o���v�G���}bY�ԏ�#�L��}��oh
v����/� ��jL/��Ʃ1�������u"�[vu)�N3�r�[v�(�=�m����"`V;���Wq͆=��4t���!v��nG��4$)���t7��+�<�����e�3�_TC�]�lC��F��9 ��¨L!�����r����yz����\��^ɟw������wB@�0�E��e!��Q��j�r�p�ܓM��=�X��\�f!4w\!LU�h��
���М�~9�<�>�m����,�ޜ��&v�q0����<�%�z?_���nLE�.@��oq��v��)fu������#��r���DC3���*Z������:o�Ht4��w�����ԑ�������H�0��@�uo�ⲗ�]���ѩ 6��ȝl���y�۷�*a�L�������g� �w��Vh%�!$��X澸m;��4��lzoӉ��H�˄��c�_f�C��c�O*Y���u)�MRƸ�k�}�T�L�5��;_/�c)	��87�P|��rl����eh=LN���ҹC��&-�]�ɥ7O�w3�"G��P�_��9��R8,}��r<������9�J�a���)�MaZ��*e=�m�{a�*N����fWNY�w�̆IJ�i~κ�dr��8J��RN|[h�g��b�<���$��ᠪ��|��.\}���eo/���u2?� �, ˇ`Ɯ��M�j����,���3�4w�r3&����j�1|��-�z�����36���y��]M��a�7�&��	A�q6�j���HB`�ȓ�:C
�X��,I\6�7�r��9Z�WȒ�'z�v�^\��u��o"`m�Ϸs��k�1�F�]��vX=}�=�+>κm��De_/��;�蠆�|����� ����U�v"�M��{��N���O����N�˼|m����<�n���!���|�g���0l���OC,��� ��A��Bc��_�/�ĄLqe�����W����P�!���#�q���A��� K�\��6������ʌ��ga%D]]�,p%�C���iBHInQ������$q܈f������=O?'Yz�pf���=J����ܣ��k��%TBp7H���I����sR�@m��Ui���Ҡ2� ;�[qH�q��ע�s-����|����]�&����&0�׉#^���O�;�@G&6�)gMNL�[ǲ��3�nB@r&F�S�D�<6n��U8���!t��\������-珙��{��{�6�mz����Q%*aI�M]��z�H�\6S����deNB���~<�����<F�1��!�z�ݿ�Eb����7�ZV�Ít^?��C��j9�jM��pnV��^�aj�4h1ߵ**�O(�H���NM�������_:`^{0߳�ص]����{W^�?��%� ��y�r�XR&����E���#�/���ac	��#�v���ҭ�[N�%�:��4��u1���c
������Z�+�6���
U�3�M&[�@#�x1ɨ>�B1u�U +��������o/�a��Tk#��R�߫(m��\'*<n�1��a�Uͫ׺R�U�v}���ss�V#M�eǗ�����p*��g�g^8K�H6h뺖ꘓ[_��z����K����D�&8}����{���Ŵ��+0��Y��dFP׉��c�K���~�R��݃�u&���2��9<���(���s�ES��P���hU
��1�G���h������A�^��Sh��;�sT�������/E��~2FZ<�o$� ��?%N0?��C����883�`���J���4�m�*'>M���=����OR�$0ŭ��dh]��w����-G�|o�4�hD�C�l���Iyx��%���
���W�����٥U��/��Z�Q��tۣPwV*���ە=%B8fP��͒��^�����aPy���}ս_�����������
DG�̣J�k����Q�O�a����ه�X���Q�_��4h���"dNY��{]Mp6�wo* �������毉��2o�A�G�t3�}u�.�"��h~�8q��.Կ$6CcQƴ> �.8)~����_4wL��@1�PB�W(N���ؗv]HY�#Vgg�Qi�:U����p)#�5փ�w���AhD!�m�ӍUBM��XV��>�zd,5��ǥܯ�GR�Ł�k&��+���|�lZ�/�g8�����3���i�ݱA˨�N�y���1�F��mz<e��?J�j{��ƛ��ۛ�63��+/�������vk+i�Q�gʽK�8�p��L����f/r�j	G����o5�]��B2�w�J�u^�B����M��V	���jk:�n�J��$����[E��5]�A�`��;��[��,h��n���Bp��ww����4��c�}�k���j�Y��5�b��R�M,p�����J�5`��HC��c�m�������z!0X����˄!�t@t��4w��l�w����_���}�`r6=��hH� {�C�z����V�8��G��ç�}��O����b�Z��V�l��X���!\P��jU�����A���mو��ޘ������a(y+iQ�Z)aӑ3,�h��iG���a9�x@fX�L��S��Sig?�Εj�?C�K\Fҫer|�{��Ut�^��⻄HJ���gg�c|w�^���i2s���p����o�o����H�ќ�=�ӢR(e�b"��R�`)�+���:3c��8����i�0U��MR�����m�7#Θ�u��mG7WP�����J����n6;!�v;��fO1Ҧ�Z�!�eBYw�*�yR���_f�3���$�Z��Eԉd���Qr�EE[�������3'L�-F\�����y��Sd��ű��lpU��"uIת$�x�2�L�H*�*տ5��!�b�j�B1t���<�8����žƁ#�sr������F����Dm�ۗ��8�+7�	�i��7�M���3�����[���8�w>��X��VT�����O`��$�ʯ*2	��9K�(�ԑ|Tv�/1�[ܯ���39�HW���Ug��t�;�5ޒ<;dM����jx��	��I9DdŘ@4"���)cE����F��!��cK<�29���W��~aY�����^�>	9V���bd���vǁO�kr5{g2j��0�.F"�vX��Aq_��M�^c��>?uTu)v��b�i\9o�J��sK��}	��U������?{Џ�>��Jg�J2�,��pSt���`_ �)�Y�<���I��f�3h�����T�?*���og�^�1]>8�o����a9�����8��+=w@��}}j������b`������ �'.EII2��z�@���rߩؼB�7���8�v��?��-p��G���.�|!����g���~'F��PP7����5�$/"i4ؽ
ǸIlu���"�@2��`��<�\��&���V��M�I�lG���!�&Q���#���{�n�3�X��՗Nd�c8�E���h��A�ktd��rX?(�7�H�SǯO޹yL���+��[��ؠ�?�Ε�i�ԲV��P�Y�]D(� �t�D����?uąwlg��z�v�������m3�@�,��������{���;�'+�OV_�8PT�ʣ����4D��mƚ�=\D����P��|A�aI	�R3���K�������ނ�� ���OLW����Sj!V���D>B�Dh
/�k�*AG~���%�Z��Ƌ�]�W��!�v�Ub>����cv=�׍+	ϲP[]��;\��n�D۩��K�f��9�Ư(�wt���M�����V��I�=P�~#F�4^̊=���v�f^�����V�<��!�&��~SRp ���͵[3#Ӵ�1��˹�^���(\���m>r�eϔ��e��-]Yɩ�W�@���x�P�)�ʘ�ɫtk�*e5��ڿ`` ���D	�%��({^E�2��>T%���w��>|�2�c�\��\��B��rð��0���s'ȕ�� ��M�n6�z!D+�L�F:���)�򈵙M��dGc�H��tS�h�>���8�?#�w:�����r �>,�����;%h��r'>�a$]�	�2b��I�#=a)z�E��t��Sx���e�� �P[ĵ�'�s��壧���@)���_�6;A`�i���X�yF�:��h�B��F��Ը885�]>=;�_S�Q�$�SH ��ӓ����e��B�?0�/�9dw�ZX����Q��k���������w�GnM9���a"���&�D��~���ٓ�rX���N�ڽ�W1�]�+��/׻���[� TXfh^���}����Kd��yw�i-��$)�_�A���
ϑR��H/SX!��-T��.�(�Ȕ��Y����1���v��$eD�9��Jd�F��"�����
����Y��g�xkaܰ'&F>԰�Ɗ�	�i?����Rќ�䰬�@Rv�K���9윑V&o�	�)D�T��o~C)+��*�ؗ%�k��������N��(���Sa��q��������h���9�H�?��cO�Ԩ-.�~C��	)���&�j�U�\��Ƒ ]��_Cdڕ��r�e�d�v��$�Dľ�*:<��)�F$�P��f*p�m���ͣ0�d�I��24�)������b ���Խ������N��FiiKo�G���*�������]ˑ��o_���r�y�I>nB����|�,�@FZ��ߎ���^�9K63��]����C$����&�{�׉z���2<�;�([�!%��,_��֓�a�,�8��%� �c+A�N�J�XYV����8#�ytA�%�d�?��� ��K[��KG���}{��/#~�Ga�J�B5F�?f�}���X�� �K�%n7�Ύ�ON�N ���ņ#nN�VDƖ�V��·>k��wy_�z����ƿ��Ķ(ɋ0�I��PH�K5���3�g�F�KI�u̧�Ί�{1��_E�_-��=�Js=�;�F��Rm���-a;�N�!��6��G�-�蔄S��2.>�� ��P��gR�,�ʏ��� e��)��j�>�'�9*����ݭ:^7>���rz���]d�J�7���m,t�B���QP�AX1�,�E��?W����Ϟ�1�a7����Ej�h�$rKWNY���b���2�D���*X���&�$��p'$r����8`�iG���1G��v�{_U�Gs��d�ł�
��F��	ë�K����H�G�n���5��ЗAM]�Ƒ	��M�����d](�d��ǹ��B'����Vv`�������ݶ�:�9��9�̟:��\�rmaE�>�� ����>��3pF}0�ǂL�Q�К��� ����u=;qo--v�$��ݢu^�U������/���jk�s�EiD�j�,7Z�w����/�rJ'T �N�F�#}�~��|������r�� �0�A�r�����=l��/N�V�1�p�m�e^;$$�}n�EF�Ӂ%��Lu8|��F2�;�o�S��Pҭj�e�`�R`�5w���(�h���VCAZ��u��=��{G��|v�ʌ�ULƨ"�楂�@IJѠ��^��WZ'Rl�~�l�`��s������`&�	�eUn�<lagndtƂC�n��XB�O��'��9��ZMO��1MĊ�|s<	�كө�ܧ����Өo�P�(�uJ�DЏ�_ll<TΓ1	Pd=͸�dn�0��,���Gw�{�MO�]�䬩���/��*C�y,!�=U���]N�9n�>r��i��9�1���m�s�5��+!���P(��"�Y�,�X�麭��{��*8���^l�^\�NH����.��(�O��� ���y��l��Rdco��_�z{�8�$�x��Z�䛛��}�u-�H��7g���tk.NXRQ�\��"���B�ph���8В��}�w�!���ዕ�䯊L9P;�Ǘ�	�횅7Y�Ɲ9��0�/�Q����I]D	{	7e��@�-J��~�5��1@�̛�/\K�n��Q!'�]�S]n)�)���x!�ɭZ��:}.V	����P3�W��/�&?2��P�GWBk�E��YoY��4!X�OR�1��ӕ���z}(�Y$p�m6t����e$��f���;��
���v�����}����@�����oבX�s��}d�a�0K_��ډ�J?�e�0�Nb�.�4�ho�>���È���f���(���b�Ք�
���:�����Jt��-��ρy ���s/���T��M�⋻��[p.9�(��Azz����[�M��&�
mPX�r�f� X�F��Q�}�����վ��7r			"��2E>�U{��b,��yM:� .Ux��9��YM2$�_s��"� ���C=����������җJzۤ��`_"�����\·��˜�B3r�@�@�{4���"����-7M����I�HH��w�u���|�< �[����w��e���	�������ꁮs����kd%c�1�?�6����GPq	u�҈O2\x��1��ݤPV�e`"jZZ'��"���Cϵ�$z&�����CF�r)�`^;����rc��s���5��z��N.�$`�h�!	�1�ew+F8�p�@ *3o'5Y�<���9���̡gDX��?�G&\_ǉ��}B�v�v%���G:�8ַ��%48	���ҵj��X(Ȧ����3��?8H��(��X�e:gQ�#zGB>���튁i�%���u��¼밫������C拚+׀,��< ��f�Bٿ;�/l]5B�տc�~綬���>FC�;zޱ��wsn�T��b&|.#�Ϗ�iԭ�*W�gE!bG�U�Ч  u�OL�8T��IO��&Ծ$���[qƸ��A*��Œ��46�A�އQ�'a���3`��涊"!
<y�p�Y���5XA-k{O���^���Bh��`�Y��|�1A�R!JPFL���Pg����Z�\I�O%<�w"U�_��,�T�z��h�c,���1n�����Q���%�׋7�kҳ23�`	i<����y�ڊQɡ"S��G�<(:Zgs'i��܍*��/oR�;9�*CSRR����e��.A�CaΙ�>
��7�Y���5(	i��ߩ]Y��|�����`���a���s�k���{�?E���(xi�H$>Tb��\<��o_4��E1��N�	P?XX�[*8\]^�\�����>�B��Sˢ������gv��n��v�����gh���.�\�{���G7�r�چp[F۰�B��P�b�,�� )�e;Uj:M�g%S�m�<oa;�G�4f��20MΑ�e�B䀞�T�e,����^�Q=w>A�ڍ��4!q�j�S�����ع�T%bR�cو��[ɡ:��7mQ8��0�wL0�s�4���ӂ^Evx����(��1��cc5)��>�h�E��������XtW[���sq�i�t��sUX�Q��%�7��>��Lz�_�� ��V�#t�c�,�>8��K��OϹ�p| t^������M�`!,6�pW�u����0TP�G�����D�z��AoXK��	��/k(����g�CCY�k����������%���n����-�v�4�}Bϻƹ�dkbk�}�.V�H�Z\b���R/{~�xf���9��~��ߖQc��5��-�a���]#։���-�	���|z�'$�	`�F�`1/�� 7��ה-�`��y.�V����)ww�b́�
���77P�������7K|t�]��o�zw�	C�aį�T��Q^�mG4&����)O��
ؙ���n>�ZF�)�"���#��"�YK��H������q���Vo;���|^"�����&n�}A<3u�&�W���s�0��O#|֤LC�ת�+����ᩢ{8�,�h�B������k����I�,��4�e��O�k����1G�q ����>G�a�e��9d�^��,"dPF����x����* i��-�U��ϚG��d���>`�s���-{�|�;#��&��v�q������Ǘh�}��?���S��*Ij�c����68���:��2�l<c��H	*eH��M^jF6�B~�S�h��Ȇ
��ÐJ˟y�Ȍ��]��t��P0�E�A�)>��>�|����M�s����a �Jf�SS�2��0r���R�m���������U�M�80\b���R0kI����v<��Z0��Q)�DTb��|Ӟ-��q`'z������K9!^��HS��]���\����u��=Ԧ�m}�d�F�4���O� r���x���C!2�����PE�W�}�{��[U����A!�(�o�]�U���_trfӒSp���ӯ-"�.�|/�M ���g�oU���#!b�o$>�9�H�ʃ� FH%Vv�(*lTLt�Qx��p�̑R�»eoΒ�(��K0Rb@z^p/U��/)��� �&6v���.F���jwܮ�������&�ߋ��+�G���q���i��D�H�jg�"�ݵL(J�y�f�	�捁iP�k}���H�]�4�9K�H�K�����h����AK�BB�o�_k��4�YR����ޒ��
ض}밐E�б�d�>mxܣ)$��!�7���+/�K@���a�NJ��:0m98Ybk�bD�ݹM0�<����s�R�yzϓf�]Z�,]�nLaF�Sc|�M�%o��*x��7�P�y���,��3�<�6�}���tT�P�����'����p�I��Tf{��-� Ng�8thL$��JKϒ��Z��ן��^���O�ĕ�g<k�OYǼ7+]/O/��ڕX�M� "�A���[l�a��<���DD����\<c�&�bCW��Ba�D�L�M�P�v���d��%S�$IB��[ʕZ���f9����y:�g�o���|"�-C�Bh�R�p��n��{��(�4��Q,ۓ��¨��M���E	E<b��+5��Y#��<��1�]�#���ؗ+�ܢb*�@ �mݬ�\�P:�$$ų��&�s�؋�W�_6Ŀ1dQ�>!}�!�G���F�s��̮���;،a�|��x��l�Rw�z�����ʘ_|��b��/���ac���ŷ�'�^�+�S�p4���D=�v�Ϙ�Sk���?w�G.T��9"O*K�n�)luc<<k(*K_��O��;����M�W��.�p4�I��k�H��m�uK5��z�l��#����qc�8xx"4��+�s��0�y0Ej�Vi��2��d�C�7�4�.c�j�^R�Z/吉�^P�(�[)+gbŎQQ��덛&G۠5��8�0b�3_����sޥفChH-ow��9�E[K��4Z�f��'ՂN[x"%��
T�7��͸�ɦ]��1�8]���#@���&P?�k�� G��Z��;���U�J[|RX�|���0F� �I�`!t���]=���
?�x��D�T����W���Q�Y�t�W�=0�W?��w��d��'�?l~�'�)5_;�yY�L�׌�pC>�&��j����M���+�é�ħ����,s���p00���`	�ۜ?�:��zd�����t�X}�i5�ג�����J��8:6���%əibl$�+�J"[8��l���zǂ��@`�k�i��r�pU��;]�Kx�o�=�!�e�Φ�m��q���J��*� �g�D:��]߼"�D���� Z�[3�-��3^"Q���j�h5t�A=�!�m�k�{�RG������6�.s@$7.[�w��S�z��}��|��Y��/_�F�<Be��s���C���_>��AM��U�P%U[� ��.�2�,$�0?�'�y`;]Fv��7X��Yc�♔0:6�Z��*���`���ޱSex���|��u#��Y�a嗮A��b�	�Ծa^�����Gt��(£�ׄo}/��'R�>�Ղ�~~LҘ"�m�U;��D�}}r

�����F��9GGmٓC.���e �I�v]�5n�j����hS[C���=��s�ae��{��m�����ύ��_�>(	GeJ ��������{AG'��"�,H�4��s��ˡT�U��l�m�:�gK�	)P���j_��F'��Y�K��)=��UV����9#g0,�S,�m��$�����P:Aj�1�M�Vް�0���) Ş��v�\Jr<Ӟ�J/Qޞ��NL�_n���O�%YR���	��\Q���{o�,�~�I�z2�3���ٙg��)ŀj��h��˧l��~��h��5�4�|m���%���u�<A�U�R�* t��	����I!�ukm�x�Mu����.#�-��d��9/5�јË\82�}���}�oc�?��`��q�A�,/��qM�~��~G�wGP�<�b���jN ]���"c�f����FJʟ㐌R=��It4�?v��:kԩ="�3�E �d_�E��Vզ3fQ 0m��P����->�:�;,��a�nO���P�,�"�>��h2K^&:zW��) @��D����8i�$��L�=��&,)�^�#�z=��Mb�_P��J����4s=-�q�nYg���.�q�"�d�>���Ofɚ���NXZ-f&������q�-]��*��JV���2�~�M���>����ќ[E�˾T���+��G�f	� #<���=nf���:��]t��W�Ҭ6ώ�s�j���iCsT��)T���n��,JB��Ų�m����(f$	)X�kʓd8�C���x&�����:x_G�T�3�@�|�!č�S4)�o�դi$��"�>�fog]KL[�>x���_��m�b�M�
k�E$Ƞ��}����D8�]C%n��^��@?mN c�4�&�����XZ�]��c6��x5�v�|�m��U��̋Fv%�<𤧧���=p���=�[`��Y�Y��H�������SK��Z�T,6Z,VσV�rT������|��-�w�]��MNn�N��f~ڶ�ȵ�H"8p���\t!�%U��7e=u��H�e(R�D[!�gU;�P,@g�c�?�V�)+��q[�Ӿს�pK��}K��}��T��33�i�ٛ�}�^�]���-����Ջ�I�����-��N��A8�]X�������e^�=�3���C��?\�c\���(Gy�k�z+Y���p��h���&RƧ��y�&�	F�R�
�Mއ�����ςC1*N�W�.�f-a��*������B:���#y��E����f���%-L��T2����6�=i���2��+&���.߾F�:�d�:�.�v>T�`���x(^��1�t U�w%�2�ABB�k,Q��.ټy��{�UY!�XR��\@�) �4�o&�E�5�^��ֲ��V���
��@ 8�SFS���2�S��1���zU\�>,��8L�N��.)��G&8VT#B��%IZ#Br��� �-]-"�� ��0p�X0�튅š ��i��*Rw�o#
��C/ɉ���c�h1'!]o�(:���O@�rAXc�����{���Ep�(������_�XU�*Ҍf�4�=�`0l���ߵz��/fL��j [) �5�m�0m��S�ɬDaϟ?p"�d24�ffG��j���MM`0�Y��W�v����\��P�I��P:dZG�S���N��FP���?�a��٘0�a徲�1n��#! ��;aoLr���9�mt\�a����-ER��)��6MƲ��BE\�}*.e����@�WT�%Po��g�0i��8v�+E`L����0r�bk7Q=R��q�Ϊ����
fK�)E�l���Xv9����nc�3��wP���� ݃��_� v�/�m��|�[[�
k�x���]u{�������f�H(�T�^����N`�x�����?@$���tTl,A<�-�Y�Km%+��Q�U��}�|��io�� ��	"����Lt�\}&����J ��=�t�!�H.�^k�e=e\+o��?:��~}���cZ8�v��H�m��d���,�]��	��0i�$�1� �Q��@���a��q�Ŭ��@8FZZjT���b�w_�Ae����h-4���0W���vQ
~�ϿL�,j�;�c��q;o�ޛ.��[ �*ҭ�r�%ôj�7Z�5l>7�RnM@������/!'m� �I89i[E���vwwX�>t�V��
X^!8�a���z��ș�� �����V�ֆ�{����]��`��4��g�%�y��&7� pb��~b������P�n	)\-�/�5Y�F(ԫt���I2Ǯ����yݭO��|I��A�uǁC�#`�j�$�צ7¾
���Lև�(i =�i8�z�k�rn���*����G��hqi%�Ҹ������V��Ґ��^��N
I�q,�X{`���C�_��ݹwj�Y��'�ϩ���}��O��}l��}<C�ҏ@�:�ė��O�B���'.xџrX���&n EY���P�=I+������9�w��N=�],,|o�\^:<w�����~~�U���gKӳ5c���u��{�lG2���y!d�ǫQ����0���|�����B��� ���;����>�����CˆD�p,��ᚵ5��o|ƻ����l@�݆/�u �xP����\� �7A:'-J�5�v�����g��b�j>�A��[ӂż��65E��*I��@}�i�m��l��A���B�g�΄��>��#��*S���(���5�(\�M����w�(k�1�g�Ȅ;���� ���˹�� On�yS�0i�25&� $)U�/ջ�$;;�I'�A%��'/*��0
<&0:N���<��M� ���%\係?���l���%R��'FV���JsH��$)?3õQ�&��x�����?!�6��)��}���[w�C�p]�{�DB@�����pH�"�`�/!�@�l��A�;R@A�J)@\�����4�d�+A�Z?�T��6��#k�5~׀8���Y�.��žiy�6�Pp�5h����r�59Ӯ3ݳ�wԩi���/U����$
�{>��6ZgSw�M�� �l��K3��/\	zWM���0"�_7JK�&�BVԴJOO7<��`?��i�u(XĢ�A Gj�jB=x��۶��u��i��Xpwo-ᲧhWl^Pwr"!G���63]�٭m��im�{��?wa�$��ӆ��',.GJK���ո���u��%�k��%TΏ��,9������/��aGIa6cY���4�s��7�4���Ѩ�]<�!�J�Æ���I�y��i�r�敐�ȗ����9N@y�[�����õ��@N�2[��&�/K100`Ύג���3�p7�2�"3w���]��Q� t8R<"2�8�cj��#g��J~�j��E��)��8#߄�g���p0���o�� p?5��. )�h��%`ͧ��M�)�ź��9`�P�RԄ�����	u�w� ̲]8�^����+�G&�s{2�[��<ݱ�\�${Fq�����~�����}2�Һ�z�֧��^�����أo�Ƙ4x�S�N�^P�[�`y̆�l�NW,HQ��].�lߩ���7#�J����{7�?Sr M�g��gL	�3��(%:@U��C�v�Wzʰ&��d��ܸM?ћf5)��ik���DcoJ�.��%�\�:⶝"�˅4Z-�Oc��Wꕪ��'!tT	��U3�UE��b6NA�k6̳�EOJ-i�a��X��Áx��a�Vb�i)�{�-�8�L�;��3(,X4���.�/C�9���
�*�f���էg�j~;%�P��@�V���mO"
���[U����S4H��1]��?/�q4[=��]>�)s.��
�S���9������l3���NQd�\N�\*t9�>�znE�TI�,XH&Xa�Z	��Es�u5P�i��o����W�˭{��pTL#�т���6���pSRLT����&�w�ҽ���'ћ�ݴQH���������V�s7���d%.�^5Ԥ[F��*��g}��۲����*>�PA��s�n�,�KV�L��\I���W�^_�q���S�5�T�Ҿ�I�.B�x)��9��r?�ˇ}����w�H%��枭H)]�7�L)ߨ]�]�R>7)QX#
V6t<s���ص:�$Ex ��e�>��W�s=���|_�bMC�S	7�;��t��zX6�zf���K����[c��:E�%�"U���2���m'�~A��(˖����L�9I���� �/�L�<4�Z�_Qb�\�����H&U��o�Ⱥ%𨅑�>&�?b.��:����t�T�@^,,�`W&� Q��õt��#D�は(ښ��t;i��a��ܨ���d� ����c�^�u.� �����$p��X�(��- �"C�kΒ:ٖ![!U�����5V$2r��+��L=;�q`��PN�a���� )����hSc� g���f��9^g<����w����.Y��	�ii��1�1�޵��T�������}_*�tz�l���2���|Mv��0�]9�\�$lq�j�l�M��9[^w�?�	��΄r,+�{�O�Q#s��Q�CV�p�8��X�t=2�s���щ���C��1�?8C��X�k,E�|�A���y���`m���c{0jY�������n��v�1	��������NIiC��:�OQS�<�XXi����[���WuK�O/o�վ{����C�;����J��wX���L��95���X�:� '��|]j��g��/��x�cNc7q4� 2ݗ;��G��(I�v<�0��p�~���]n�Ԯ92�g�=ԝ��q��<���^�^�<$�{����j݆tD��=���F���;�М���Ɠ��9(®�e����=��6�;��}C��c:e!RE��������3�>-���<2��c}"�
��B ��@g<[f�8T�`X`��}���|�<���Ɇ]=��2B�ֿ2��	J�m��{2�J�iw���W�_<�%̰HMK��OgT���\�����c�Rw�uۮW�j��Ǜ�VG���>���ͺ=��W�D��ڟ�ٴ�+�$r��=��3���*���~- ��m��v�p�N�qq>�B��F�����y���g��������p�����訜�ONn�veA��̒�A��tp����]�ө+~`O%���3㤺+�iB0��ɠE����)�fV��Q� 
��d2=�>�@�h"ѠF�i�;����[�)w5�u��>�dC'��8�P#!���(]�>��]E�+q�S���B�D�/�h��i	+OK�V�
�����%��A.Λ� �p3BQ�sB8����U�.�XP�AK��ݰ@L%�w�:�ۥ�P-�T�P��u�ua���9.h�|n�"�@2�n�;6^��~��Tg�x�s�e����{��|��5��e�k/^�(�vƼ�f>/)��@��%gެ�O����KǋV��8o��5���3s��%�=g�0�_����6�L-B�V�2����G׈&��!��^��W-
��`�3A�~4���c�y�n yױB�����F�k�N�E�"�=6�C[�3ka�n��Z/+�����q�L#�;ݸ6�^��	��b�F1��9/�EyS��?U2p�|@�D_ɡ�a���Ά�5�\��Փ*$��V���t�@�8���g.d�B��LQ�ޟ4o����[�F�ԩ7q@�����j����pP�F�������1B����#wcD�If��ڃn�L����_��y�~���� ovU�r�x6:N�0?�zxL��Z�&���<h�n	�O;�PjT�(�at�����p�)�!����͏Fm�d���?�V���� �+��NP9*j#vI.�[`b��k�Չ*V�;V��ZUU�=S=6�d�w-�]�&��s���b��>X,���&~�$v�*�=L�Cl1��{�޵G,�˾,��2#o���6������=��x�8��g�7�Ҡ����V�v}`����ԗ�=^�#���'�BaPt�r�����Q��ɐji��r@@���]��<�J�<I�`mzI"�횅��tn~��*����rѠ~B2D��ˈ&����)[�=m�U��2$/�B;v���K~��zA?R���ѷC��4E��%A��{P��%癘x�͢�e+�Yɦ�~N�M�q����"t�Ӈn�3z�g�o�a�ߙ~����	�*�ܑI˦4��R%�h(A������K��1�J�NWz��hS�LZ6Ƙ�i|5�cԳx_d�/V@O�Y��ɘ�#D�k6��!�;z����k�#n���k���]���o*��ќ!
���rqR�R���:]w�T���1��m��ϼ�z�T�q��r�8�B!��ݘ�5�� �L��U��B`�R���?|w��*4�.�g����U�C�o/c��+��b��vS�u e8T�C�
�^�$:��4�l�4��BC��
��est(����)�9N�2|���͟]DM�2��E)k!�*��e�C�q����*��H�_:�="���/u��z�<��'�~���֜V6��������~��o
��'�Y�+V7:n�i�Č�`\���-ҫv���x �6�Uy��8��Q?BèH�ͮ'Jף����[���D���N!��:�2\$b��W�$	�8:D�՘����\���Ǟp��S����^|�f�j1a����T��p����)������ܑ�\�����S��fC�{��hb��)�q�@�Eb����Tq�w�n��q��
����l�ZjO���'nR�jOR���,jb�(zJ�HT����1�v"X�na�ң�5����׾�����rPI������F�B�pѴ���E���o�i�N\�g=Z���0�\��/�?z��ėT���ï��{
J�){���'HV1X'r`B�o���݃T竊H�����pv>OLu.�
g����xsځ~Oi8c����~�PW�d�s�z7�s��5>�i6&xwH���Yn�%�?(��P
I9
i
Q�`g^����\�M���$p��;��Z����_��OH�$5Z�Th{nt���a``�%��9�5��&����$y��s�l���TdXfO\�~������k�����fr��w�#�}�vF�ܿ�^ľ�+z_gn���n��2�5�
�_�t3��))����~����4�����W	�GW)H�u�>����0ߏ�d,�	8���s��`h��TB4�,UL�|%)�ܻ�wZ���̭?��?l�>C��W6-����`��V|X��g⺨]�WG�q/4��M���r� ��i����bbu-�L}s��I竿�R&�3��qFﴵ��;G<{���|�Z�n�1!�\
�Ù���e���H��A�x��/�"�����.�/da��X���t�z�jZ/�<#n�	���듬FC1��[���xJf�������KL-�!<��4��C|�"q����{r�����=���lgfk#Q��N�1ȧH/�'���W�Fl�(��!+��8w�Q�L+�������3c9����g�?ޫ���o�y�%�0ve5����r8r~���\�~��ޖ���8�t���u���V�	��u���l*���a�-�����B��0S�ʤ��\��bf����/1���z����O]�J��tR���'�lό���z�RS+N��-9�g�ːzl_������ ?!�E�z��ߜ�� �JI&�{J�V��ٹ`�.����-2�>-�)^��u�nD�����6b����L�/���4O��qߢ�5n�i髆*5����+�p2B�g��ظ�Ĥu��5V��K�yP��t�h�g��Jb qȗ�J>�$������ˣ�6�xx����T��x�[�d�AH��$�bx��Q��p��'F5�,�9R*SK��615���"@$J?�~�7_�m��.�U	�	�<7bQ�٨v$,j��iA�q�{�������r�7%�띴�uW�9fɩ�[�~�}{�"Y?�͋\�^m�܏��he��y}(?�U�R��'���E��7�a"a� }ꊰ$�����UQ>��S��h�< 4�oW�Y���B1��@:� �~��*�Z>�K����a��?�e
p�+�V̓�z�� I#I�<��E�,)�"b��|K&Y�Z���cf�ob�)𧽐��B?�h����?̃,'�e;�>�!�>'����,ݰ+�F�F������(��U��J�-�DC����+���b�nR�1���������F�q��o�o�s�лwj�����L��c���O�}�9���+Xo�]&�i�6��;@^�z����ɐi=,oޜ%?��0�b�p�晍'μ+�Ap���ipBBCh��l{��Rի����&l�I௿�6_�u=�g9<jU�����
���(���OWp����R��4��J�>	����o)�����~�txr�_>� E%�M�k�gG''�P��q�5[(�z�R���a�=E]1�ZP*������~��↪�d��K��W�|ouT�D7ݣ���G�J�y��<l�x{���9��X�P���ݴ�j|v�W&�]3~��I���%sl�|3���:��z|����3G�p�~��Vߌ�Ky3I���~gpk���睼����b�������f��)��|s�ШuD�t�4@>U�T�~��м�VR&)Q|�L݊z��A4�ʙV�7[���.Y�PI�f1�������:�͔׆GW0���@��...��/z���D�ʕ�������e�E���?LFR����*�j-�Aʛ�p�	9�Q_UԯMw�����2���!�4H7��4Hw���)%�CJKw����{�>kf�u��O�j+���_O�Q��1�����+$+�z��{0׭1Z��"6UL6��C+4�[�pf�k��&kN;�NP3J&I��"���[���lWK��i'%���G�3`V]!�]I�6����|�x�	����|�^��W���owl��m]-�̕sH�A�d���<�n�E\��#�gݾI�W��*� ���k��X��D�6��i�N.V�W�v�00�����o�����g��'P��h9(7�5�9m��.]p�9RL��ǒ�\�8��m;H}�A�{+*�F����ࣩS����N i������x_����o7��-zK�}�_��e�Վ[��g������'��lg�?4e�:����]���#S��J�x�K��GD���J�/>2!����B��4]�Rm�f*?���m�W����J!#�o`�����;S�稑�=d��������b5=�-��[��uHy�2v��9^���P8.eȧY Y�UF)E�A/;W\�엀�sI7+K;<(c,p���PFe��f����n��Dɷ�Cd6�ê&���0T��tԘݸ�������f��,��C\��*���L�����G������x-u���u5���E����Z���eȉ�b��dZd��X����K[�׏�����7L���<=�͵||�ڬ�P4��Ӂ�xMƜ;�Lղ^�T�TeMv�#(Frl�[����C�1�&W�/���������1%�I�I >��KY�m)�/]|QݐIt)F5��0��T�� !��t"SN*E�������ͻ����J?jj���H�Q0����-B
�i""#�'&�/�ܧg�����ɾ��c%�1�õ���Fh�Ъ��E!� �{��+W�����g�d�h���a��#Z��%����y���3���h����پ����C�`l�~��(�`^ 偣8v5G�_n���VY��r���kZZ~I�#!��9�ȝ襛�������?s|MB?\�����_ �9�`-h��� ����.p������*W0�V�J\��s�����{���b��-���Oҽ:�?������u_>ӽQ�d����6���p�+�OX~-VB�)Նs�;5�z�����pNc
i��������1v����y\�Ư.�b��xyE9p��Xb �c�H�t����C��Ȱrξ�ЫӶ8)i)���d�N|��)�BI^Ábj�cն�g�w �>�Vp؉���qS�ػ.�GG�����P����/A{KK?��ّ�����W�����ڥ�fK7dCU(���t��ݨ��T�j�J� ��Nɧ
׈�%����U�R�AY��=����Ӆ�k߳��ΦI����i17���y�d<��d@adL�IV�,�
�U��ה%Yia,9M�q��80ƫ��uF����G�3�.��p�7ڤ�e���a���߹�S�2s�6X�w=�&�n��H��6��E�M���pd*���|,�"�iO�ܞ�|:����3��K�?��ݝ��z�plSv�lc<��q΢�[s�U����t�DLE�Sr���5���N��_���a�?�TC�^��^����� 1�������$dFS�������[�Rԙ���6���/�ӳ�peB��=9�#�=ooe���R�櫓D�Αj#LI���"�F�~5j��+���Z��W"%"'��'+}��3>
�Rc�,�֘_�c$d����p�$���'t=�4�҉���WWD����p֢��l,�^2j�����lۨw_��P�Pz8����e)K���h��<5 U���Ov��[[[ԛo���w���u-?�}=�4u�,i�l�w	���,ư�gg�o�l ?�ؼer$���&���,w�"��b��Z�S�XQ�>T^[t�����5t-�~p�'��}I��(���̗�� D�ls�^(�*��5A�0�I?>KS<��K}hj��EpU2O��'�Ҁ�j>R�E�Y(�y�f)Q4f�Z����B��#!>��1��, �v�fYv_E��wsw�V�y��K����꒩~0� ���c�F����}R,*ɉ��N�CZ��.�.��-{w>@E���j�ÿ�X����cc�����~׶/�~�=��>�'�2	���M�_�N�x�o���ݣ��Z�Cħo���i�0��8�Vj���o�S�'��&<e��6N�!�{$��ʲ�	�y(qA)Ճ�}�|�6+Tƾo7��Ҧ9���	�JT+5�@����7+U�!33s{�����d[�T�ǟ�i���m nlM:~��ts?���_n R�@����!�j/�<�!��z�T��Y �k�]�J�&�����V�r�9j������`R�/~5ޘ$J�3��o'��۳��!UBzv4���HV�:AL�1+������P�J�gqj6�'�T��hk& UB��eQ+�M�L_Ǜr�BK*+�q:{ɻK���ל w���\�d2Wgq��9I�:Y͒����b>�:<�_L��:�����tk'G韟��$/��J˵4 ����\�(ڜ�S�IT��>q���Qе"�xEEW��S@^ ��M=��1�I?}�B�T q��rlq&F���G�+�i�q<H#�8��)v0���ߺI�J1uc���s<2C�ǴC��E\���k�2�F��JB4)ߒ%�m�~�$��f�r�$���8���JsuD8AE�1g������Ąg:�(\1��^����Ŝ�޻=���(5Z::�*�Nt�o����#"���;���M*Ypv�kW~��ܛ㶊���W�42�<�/�h��CT|�ݶ߬��b�R�1��vD�XH�1�]I�߾�r~���/BD	b�������4?p?R�9r�Z��W}����ud:�Z����٬/!-���h������P�@���1���K{F��9c�X��l:-��.f�$Es�^&j{�T�?mX�j�N@��G$7Sv�ٸHJ1gL��]�s�2(��BÁ�3�S�R��ѷ#(�+�Vf�b
{�:�i��Y{��_�&d����|�9�K�>�K�E�$7�E���l5/uS�. Y���*��Dy�7<����}3����>���=�!��I̹e�l���r9�L�?-n{�Y�������T����O1��)xBbL�>��}�C�D����L�L�^�c���-jN6J�T�,�]�'���T7Ξ�\e��%J�-X�R�0Ǎ��T6��7ʈHd�Cn��7~�u����Q��>۳�z�r���ɪ�����L�n�ʂ�#-t�#.� +ʑ���_��f���J�M�Ĕ�f|Q��m�L�Ep��%�q0Ov!,\j!8�v:�E�j����Q쀔�UG���Nhf�~ْ.�ip-�W>��*�&hC��������̃�S4���*Q"���r�E4˾��Jr��S�@��6Q��:Z�9P�d<����@�9������PjC%�����+٭�r�yI��$R��Ƕ�5�)ٸ��d���5�pK��z���<�����7c w�9���b+@�ʑS���&�����(�u&R�!NP�F.`��G%k����7�����S���'ɲ�(�Y�N+�+q�R����_�O���l�������i����oy��C�M�/ɴ�[6���;ļ�c���}$�*��hGAޤ���P�1�0- U��w����%eS]�6��9�m#Aw �h.���ٟ�H���r�ma���H/`��iɊ=�0��N?쥮�f��P�\k?�����5��`�����M�/���;!ٴ���C*�ɔ��!�g;�m��62�D���PUZrlzY�X���D^m�ԛS� S1V��GA���<x7gh����᎒�X�r R5����#٢�לn:�s��0�y%�?�XG��=7���ev@�VG��#����>����(:�5�����X�v?R_ k�> �.W@��S���}�������x�%\G5�ŞpN��Q
!e���r�*���[��e���X�`�H�3h��d�7����Å1��a��h�s�����}rA��	���闫m�(��K��>�!��:r�P������*�cAj����NVe���/6��s�b�tp�S�+)úm������5��(�v�>�q��h2�)������6+�G(�CmtNLÌ���ST<�
nv�4E)��M���X2��)����W���Y�'a�v4�QKAʟ�B9������|�_��B\8�=���G��\�3�t����?�5;�"���=�Je߬�>*[����*�~!��d�iW�/��䉂ꡯ�kpu*жUn%��"4����y-��*f���y���?�e����Ю�m�)�u�����]���7Ek�x9!��w���Q��Dp�lu���R�~��t*��S��^�����q����=uM��!��֟���ٔ:(C��
$]�qM-��3s���@5��X C������?j1�;���騪�7��Ľ�`��B�>��'/V�(��lt�J��+0N+L\�5�o�|3^j?8��������D"�חxA�����#���D�(�ϥ��]8���7݆�ُ@�~Tѻ�_<y�hz[�/0(.ܻ0a��˔K=������_n�}�WQ�GG߫&�����{�{��WV�˚�始gm"Ɯ��8WT���e�\hMG�*�alۜG�ޝr1�%;(e�Lj��5�l��>�k�>��1I��P�ժ�@�s�S������BZ\뢑:2�����e�L�[*,LL�]QC�kq�b'q�E������w�l��K���cvj*�6
�{;9�H?��Ek�7���%2+^�)�7���+V������g&,*�X���$� �y۶�qB���$���M�z��0�ğ9���Wtl�+��c|�Nڟ;1�����w��e��g3X�d��?!��;.�������|fb(}�_$���}Zx��E-��`�W���y��z�F$�Uhya��a[��a�tqŁ%�;���Ā�+��b�^it���#�z��y[)��AR+�~�y^�z�&���O������i}]�ꎙ1d좊��o~�;��o=�s�b������(@J��t\{P_���X;��FXW1��b�����7�3�õ؞��������%NV�1jj3�V�4�C��;�Gg՜��[��B�l��ը-TL���;��Ɯ
����c�6|4ىLL��?ե�*�M�W����-�߃c�FH��%������(�Y�ٹ��R�lm�ف*	*�ѬY�jw(�Z�+����dO#t��K�ۑ���a�^H�+��YZ5dΐ���/�=<�Ck�nLpM�;�#��ɥ�b�6���k�[������㘺E��R��Dگ�mt��$�����Y�f�v�Y�r��@C��_+�����)+}C�˾Є��s��5�$m����9����7�@�rR�ί|�����eX��]��3+���M(�c@f�ݼ��QQ��d���p��)�:�{�g�O�ŗ<��$�H���xE�˘LU�]`�/o-����
r�ZS��\�B���z�Ĵ��K�Wf��kr)�o�1�+L<��/��k(��?�㪡٩8mV�>�T���X;�+���f��dߌ&��N١j-DU�'G�V���y������*/�ϔ>���-͙N�=bM�X������8�8 	B�##��l�dy�)�r�@MM"�>���8���~�,���X的�3�|����d͂`A3c�Zq
m�$//���d��xB����Fy�!P�*F�WGR̔�:��b>�1�ݕvK�4k!��zˑ���k_{g�@m�$e����w#_���_lB�E���,yfJL�Z�y�zv~5E�l���1��b�<�jQ9<Z�b�3L�����{� E�)� I������B�y\�g�Y<���FC�K�����v ����D��k�%��!��Ѷ��
-S;���{vӹ�*t7�XH=]6�Ƙ��lU�^�Q:�	��	g��,$6��v%�6��0��������ٹ��r�c���^�PR�m��}�n�i�)�H
n	}7�r)�_����8���m�n�J�>$�ܕ�u|��v�e��_dR�<�?zp�%��(�ti�-/F�QCY�5ut�M&afG+Y�w��k*ڂ� R�0���2��5qi>;���>G{.jA���D�bOܭ$Y���a�(g�����oW�^A�#�ӗ���1�$�'Λ��EY�z�������V�%)��-���4M�)�{DH����%�6�X� �T�!B��[���2-����V�
on���Pd��dߣ�t8ymW����a8s���a^�j=�@�i��S��Ƚ��T,
��t�������}#a�g:�������'g�IN^a�\;�=��~�t��4R����y�P��pbӵ�����F�cSsmR�p"���}Wu����� �N��]ՙ������=h����t�R����ΪIڌ{`�������*N��YU^���u#�5�X�o�&(!V~ Ub,f�7`y�o���SA���Y8����]`��`p�>���G����(��Jd-�\�:�#~��  %5Osr�����#9{�S`��}���;q\Ke�k���� 9}�5R��>�C�����9qq�xFAB=TP��3����#!#�\���5x����Hz|���)5�葽ڞs�ݾ�� ����W�$�q�o�5|w���<���$�Y��z���[�s7p�@�}���\X@���a���Nzu�lP���מN0�akd�� ��.Y����i���|b������������/o�N��I�L�,h9➼q���.פ�~+3�a���@�a;�```|;��.}�N�*a	Dd�HCh5jp�����j�u�|�	&>!QQ��Хl�xA��T��@]����u���u�J�Q%i��b0��~3(d�D�k�/�w��Cx+�4970L�uv�|F��_C�@I���&�T��	iv���M��h�%�Ѹ�ǒTa6E�>��?���e:_|Wy�z/��R�P���E!��6
W^������	E���c$+�� ��p����,~ުi;,B��Ф�>PD�*`�������Pf?~Zf!�[��}�f�t|���T���v����$#eJ�I�ß�ʳ�z%��Q*-Ǉ��xֲ���@G� v-�t��:>~�0�W�$�Ye�啙Ժ���ƄPY2�b��j��4e{�Y~�Cɝ�i�.$S<���
0l2]��j?��[>kY�S$$/����T��\:�x����64�=c&j/��^(ŖcV�����&?��-�Onm����*`�������s���<b����Iu��B�g�R��l����s|*WL�炚��/FE�����d�c@�d�P���`��T���)g���
߯���8!k%�w��7o�F!��"����X�|�jI��?�l54R���?�Ly���,ν;��L�9\����{GRV��a�0ZC�!��,{t�w��#G�*P1Ce��/)M�s�F$Ǆ��b�a����P��wpv8h4�@� �G��T�T���qlJ����7�` ]�4�P ����x{��7�o��>x*9��Mڍ V�wn��pOG��P��d��:�tJ�L
�\b�M�Q�O������%�:d��x���Ng��B��fưس�����P����\
�$���'��LN�}�dj�UA�J�����1�Q[�����7D�z���d���5f5�6bQ}�fuK��$Cg#+lQN�L+��;�y�r�]��
�!}�}��8��}���0�K1�Zlgs�\\pˢl�ptNLNn�S���C�N�Y�tݷ�=y7r�����S0�M���Mw�m̃(IX����Z&��rgg�\����H�����ڭ4��2>f�U�wW��Ѥ�j��]����N����Q설Il����-���'����ԅ�H�ԧ�C���=a��>���>����[9�LrP)�.���� ��E� �$r�t� �gZVpӔ���R'ڹ�{*eBe�gz|�x��C#��b���儠�p}C��[��l�<c� E/XQ������]H��2��G�ȠZ��뤠�a"���j�ÉOh��l��2�_W�GJj|�����ZMyM]�=F��}I�{
	Yn�I�����U������������SI�5�#�H�>���OG6	ۅ4�]��FT������6��0e}"�)����{~@BBZ�qs���A����j#:��Y�?֣_���_��ҕ�wm�I�<� me�i�4-J�M�Cao�v�� ����qUZƪ=s��Z�L[n2[��<����,c�9D_M��9
 �� �too2�v��y6btϝ&h[X]A���cPP�b��A�kt �6�䋻
�G���E���z����x灝Z��R�	ԛZ�Qtǭhgy�N^]���=I*$PZ[X|Q���J=��Vke哲]�[V.�X��׬�}��v�U�C��((�dc?N�����B���\�SU���Խ���oJ/$�F��+-㝩��>@6�����e�ZCMӷ#6��b��C����/�V�4?y/^�|�W2e����g�8�g6Y��f�ن�r���X%l`ɱ�|��|��:\��Rh냉�!�����x��S�����D�!�=�Hn;����<�JZ���>�5Xݽ��Ë�4j�2��S	���ﾜ�'����p<J����H=�l��E�`uMAe���9��DCC^l���3�*�з��sH�ܕ�V�HгpLLɯV{�F��1���c��	DK�;�5�䡅��h:�k{�ݾqD�kk���r�g�a8�0��y\���i���$����#��(��Z�4*���[��i�"<oY��֝b������UT^ �q{nx?wJ�b��o��KX��B��	��F��!I�
��N����<t?S��Ǟi��)�{�m���屇ʴV��X��3bDDz�Kt윟�A:�=��	�a�|;o=�c���0#*��S��n	]̂Z��٭"NyA)�R�V��l#��j0w$Mns��*財\�{ �~��v��bÞja����:V���9�&(�x�V<��̩d���0�=�4��-O�}KH&
4MlY���D@����j[!�Z`'��z��lI���)�V@�c��-.A�h@rh#8���I�?L�"�ә��ȉjN���*�t$�ou�@$�E���!h[ڧ��敧��Uy�[6��f=��,�[��ddd��܌;��lG��>����3I��q?�a|�꺦���߮�dmf~�}�	�z{�{n4��n��jo!a���$s��hг�e�BM��m͢�����
���4v�l���*۪�vHH��U��|in~�*�$O��d/���6Τ��������s�QQ�(C�R]��e�I��m�t��(�p�>��{^>����5�}�#��i����S�����̳�N�A��{�5����{�_�+�K"jn��a}�'�> �%�	�����=�o���:�۞��)�ʫ+�Z�p�T���.� �σ|
�m�w�̌3�oP��I�3}~�o���M�eF�Ma6_����B�uu��)s�+�}z}r�nDDDhz[NA��E����J˲ܵ���'Y�ߖ��8Q�Z�K��ba�B]|�IM#��ݸ��BU�1�����  �a;Rw���w�8�K���ܬ1-�Dk��ы��tɫq�qw�� �����󡈛��R�?NH8�R��}t��7j����}ybz��` c�S�Oqss���қtˤJW�L~��HMG���a�T�2~�����n�2�#o���Ь	��T|��^���Q.R��;R�I_	qhۢ�	7!�O�Iij[�:m��"0v�w"�ƍ���#	t�����b��qq�x;�vIcpdC7B˒��X�,M��bQ�1E��!�	��"���-�R;�X{G��-,�ãX��_Rx�� o\G��X<��V!�K:<����+,��E1m{i��^}x��G'&0�5rK@��<�@m5#�z&C�z�k���/q?���-~�]x�u�?�����4�͑Ğn�G��6�S��=_
\*ݾ�3S?oOO��X�ŷ0Q��+��H~}�hС�O���!��|�ŋ�[D�0d�Bn���i��a #�+�����L� q�A|�:�g,͚\���TWW@��iO'����%�O� @FY�Q�����.�d���3�}��sԘ�XPF��+����9������^U]��W��G_<��;�3S�_�8�x�	�'�/T�º���ALŽ��;,A��r�'㇀m��L"����<�����;�_a�b���t`mS
#��2:�p/�+�c�;��}_�s6��M�+2�XmE�;=���w6�V�<�L`f!�*D�d��;)�.�+lG������0����m4v�f��4��|)���ìI��M���1�RS�C�fa^U���d�N"T)��[��%TWo� g �]h�I�bNUy���npٔ�W	R�>[Xܝ����qe 
�"?�"%�i��.sc�0�@{y�g�P��ѨaaE?��� ��/6-��tpB�(���Z���!��8F�'_���QE,�T����J��ʌ��Ṱ8��ZFFIhtЏ��*����a/��UAze�(Vx~F}F˲�LJ���<=��.��*�u'�E%
*+�0�|��LX2Y���������2D�=C.����h�v6�ح��FK�s����B���6��N��.+7�a����Kr	z�\^1G�B�ק����� +ӑ�}i��{x���ⓗ���8$�a:��S)�m�g.n;��b�@�C�R����7է�1WK1�Q�&`v��
�Ջ����XH)�2�y�-��;��zX�C�-�&�)�-�u�) �r.�o��}�Ax��;E�
�j�J��Ŏa�-U��*��pmc�eo�9b�P�eȃ��Qa�*NV��.���'8Ip�#��@6����`���%ǎ�y��~��E&�#�vb��(!�F '۶8��N�+`q��7U�P�w�*_S�]XP%A�l��m$>��nC���?575�4�ƅY�zG���U�)⼃z�q��?^�S-�&ފf��\s�y~�������!�G��c��v�B�Y3�h)pQ%�m�7��u,��c�X�1�����1�u���T��#�f[�B��@G��G�sx�����(W�q嗻�+��Sco���`�cr�������Z폴��f�h��*�?�z?�%�?M�4��я�"
� p�vs������.���}��l3.�{n&��xM�o� ��j�O�To(�������f�%s"Uۮ�C��A��^N�~? ���{ʒ��)��Q̯�̋����G�j~/E�����L"�_��*���9��������6z{�:Y�L�CN�3䬷�������"i��g'ۼ���g'���߯�
��Vݶ�D�a=�QE�3ʇ��	��f����j�Q��O0M�4�������U���C�a�R
o�/KS7/��xO�g���a�p�B����F��7��0���W�d���TU�^���)����S�#�⭟��A�5�5�&���y?F�^2%�q9��`T�Xj�0p�T�6�����8���՗��4.U���6�֣�>���4��j��2l,1Ҭ��Ƭx��T�AC�/�
`[~R�A�M�0�W�΄�ቩ)�`�}\�B����/����;B��q����}!����S<�d=��_m2Ϫ���q�}'^@I9�Ŀ|�$s��*�����y%��Qi����?��������V�5�% "(Lۊ�6'8�ഁ�X^����'v��Z\G�m�oj�QEV�R|�WiD?��� ����E-  vP8+;"]�[��'��2(�k@�z�`�m�gN���;W��^�B�~���3�@ҁV
��6�Ye�V�|���	���2�)r������f��ܧ��]��OĽ�7C�KE�N7���~1=<�����К�06�����0ڍӼ7<�dQ��E���333��Qn���ө��ub�=2G�*O�f�|�>D���>$��0G�m̭դ�d̳i�n�W�L)����l�Q���8B�>Y��׭V��wxc����p/�=���	f ]:벓����������	S�Y ��b���Cn�c7�rf7c�����wiB��nGYQv:�%P���k|�籮}3i�2���]����O�Q�%��N+��T$$�ǋ�����K+��RP�*(Ϛ�ʇ�oE{�v6�� ��e��M�cV|>5*�����]!?j�#~�vD�Z��g�d�Y�������{�䱈�f{��u�D.���Po�����̝�ǩ������/M��bCP�=ܬ6<P}������z�S��$���eHr��m(v�ZH�;�p"�P��|�_��i�祢Nɘo�v�vQ�0[O1��dB}�,�=2_%�Z�I���Exp{Ǵ��Xr�?�n����?蹀�	�z�䒵5�S�h+�&H蒅m�B��"P��\;��bT�w?�����o�@�e=������B�r$'�����\�w|[���J0G]w)!Ww4�1�^�ȔzT�w:���63��4�5����k��,��������ä�M�f\:O�(�A)� �l�F���m��K�kl�lѻ�!j1X4�����y����f����u;ۆ	���7cC��M��`���y$sP����$�}��-<������
JީDZ4�L��
���22(�*vjM��[l&`x���t�9��R�o���H���WS�~/)��#et��Y�I$�p�H��i�X~ɽ>%<���s�p^������7F�'`B�R�+L9�]@-�EQO�F��L9�gÀ�Ցߡxj�7�1<Nl�Q��"ʥ� .�Vy%Ιw�y,��<d+YT~��S���|x�9��� ����@����w��w��_�#im�G^���Z	�"�ԕ�ѕ9�-��L���o��A n0�`���E�Y'�瀠��-��������;����ӱ����+j�f�!��]�գ�t�F�c�jֿ&�c�6,;���qvv������Vr�����&,�%������fѣ� /M�ɢL�'����&i�\Ϸ�����%�
��`	k
��0~j�3�qh07)
S�>�e}
ѱ0���8�WK�I��B-G�Ǐ|�=$F�(|�d� E�F�I��:Ben�x�R8��x��_���o�yiMR¾Z�I_�2�j? ��;���|#"���{"��ב�F'����6v>��/b��Q���7}������h��-�*\�?��S��r�؈���Di|����W$!�ڬ��պ诌��*p9w�mn�kYgMևJ}İ���0�����H{;G��T������	=K��EʸOV��YV"P�j�OM��l:6������M�Y0$\��_pb�[V���e�U�JWO�2u3Q	b���8UІ���7�w)�d���_n	?�o"��ƈ9��*�Ud�Q�[���vB�K�e��[�S�^ÂJK�J�pG�K��i���/�q� �<�[�ġߡ�ĕ���f��*����F��c?�c������ZnRKp�fڀ-~zDG��ٵ��Q';��	x����Y�~�B���
��~�U��p_��ȿ+�T_ehy�����2�}3p��{�=�+��-UF�������R��a3�!��@�Tgg,��TtN��Jߔ�'ӷ��TZ999 �#�\��Y�k��*;��I�}�V�����R���}�(�y���p��b�C������&�CL��L"x/An�o>.B����S7;,�f���Z�=���n�B�alchh���@B�o�g6ߊ����3�cd��{��_�)(]���������GC�6�Ti��,rc���݆�u''��)I��	�y��Ĕ;u�7��#�u��k�;���X� ����_��O�Ut���5���'�(�{�}u	�3�]�8����fc���`)�A�+�|�oM����|S�\X�?mlkSMv>�t@�QB�e%a
�eF�[�4M���k�Ц��fs��p~��"q94ʒ���Ł��εX�/��-*�|�j������W�}��Im�+���5d=}�[�a����޵~[ؽ��riD�w��
B�p;U��U�߾���R��jaM�z�G��G�;�U��.[Q8�7Q��ʂc4�.���oO��M��t'�H���c�QL�?9��K�A��~~��Mh*����u�՚"/�� �h�;�1_���7�Ͻ��K���QH�:T��'��$��^��K�K�,v;�XP�,��o���T@C��;���f]Ϝ#Х5�5h������R*�Y7��S�s��O6{�����훿8!B
�������������P�����O�xS.%g��ǘ��z9�� Y���![� �|_�'�Rd~�[�B���~���VY@� >�!s,
�F"��pM�f��/�/�l:���� ����3�Z�����έ��\�I�����"`#�"�	�Q�㑠ћp�������)����>ޟ�/���n(iq�s��5X��}DTH���5�\ρ�/#z�QM�T���I*�Q/�t[���E(�-��m�yި�r��
�������G����8�
T�[�Z��E_
�GO>d�tQGwUrn�s׉���4�ĉ��N���^ eC�<���5ɢ���%�(��я�_�S>&�����9��l������~�kb���4��ΐ�Џ�"��g9��aG���a]/�"�@��Ǳ���/M�IPl���q<���r����'WW2Ɛ=+�$�cZ-W��Qy����u�;v�x`���n����ٺ=���Ģ-��$�Z�_��ZH�^��5O�`��M ��Yʥ̄*y	G����ɯӍ9���3U##�6l����w4؉.I1ə`�[v��o�?*�7�Γ�}�y�m/3T�������@ko�����oT�텀��m�� x/�AbӉN��kή�'�X�9�r+,h���b��)�aե:�wJF1	�}������0��N+��:��;��	y�% �y�7�S��Ft���;��F�7��t�VL����l�9��J� t�M�*4,h�Q����-��|�y3��VÉ��<ȼ������Y��}v���y���l����C�7T����6C�\�~0��yL��v�V���χ�8\����.+�_��.��6/�I�m����J�D���MjG��Rf@�k��}k�/�*,:��ġV|�HK�c��ɯd��F��z�Gӵ(��f3�Ԛ�}OO��j���T�J��v��{	:߈'(��ݛ�W��wJ�QX�iVw<��[�/=&�wҵ�むHw���M�e
#���8�y��x����Xὴ��Cp�i�q�$TlA=�ƄpI�*�:N����R­sXay\�����-q)�D�Q0^�p�2C��x=����^�߇Nc8�\=��XUl��C��C�� T��A�V��#u'��dK�~5?�YW�x�H�v��>Uş�l2D�v��������?B���	Y�ͪ�-��m����׾���L�����'�y���?o^R,o$�l:�,�wS��;�Y_�P@�?"ґ2h׷��>8���}ɫ�����cV^UMu�Ӈ���)n�(ļMo�x}d������Hާ
!�Ôp�m�GN�['����
)B�*��HO��/���h��NԒ	�����*s����
ֵ�GV"&Qc���/��{K�-ڵ��vКR�ϸ^�w,�o���Zu0�)��]�C��$������D̅c���h+'`$^Ƀ_�Lw[�v�D��u���d��Z�����;l��b�Έ��A��`/����%wW2��ё�(RtR[�r�b^&�@]��^x�wJN%϶�4B����k�䡡����-t��2��(LR�i	���J^��d#^J�a)��մ%�$ŷ��	BJ���⵲O�iG V��=�y����������@?K
��1��۾*��*�XZB�c���L`:��kQ�z�%3�scUKk��';����RrGwX_��1�Oo�i;��Լ�F�Z�a��7�)ߣ�(FmQ��D�Н�  (��re��KN��/��;:����:U��0��}7�;�R�`/@��;��W�Eӹ#��3V��ٖD��͆qn�����SR	C���R)�����$���j�O�ɍ�n_�;� ^?�J��'���vޛ��O����݃�oN?�����1�d��K+�ؗ*�/��$\��o_��-�-��0*$����~h����־���(���|D �L�eP�Q׮q(����nER4P��ݝb�݊/����N��C��}�9���L&3{����~��Z��q1@�%�mǏ�|`�`?#ֱ��Tr�NH�Yg��D��e��@�_,߰ƙ����� %�.6�ר������P2��8���h���m.� ,_�S��M�\�fcX�Qh OK�9�-�0�ߐ_�S��x>�y�F́{!O�<5�)��[���f��Q�~t:��"O������K��CŚ�޿9��h���C]�c�m{�l����_f�b	%�MiM��y��G��WP�����O�v͝�.�4F��n~ ���8��)Н�e�%E֙k�*A�W�/�����ًYM��j2���\�L>��M�|nf��_	�|oK��7��V�m�*�6G^o���2v���]����K�s���L��^�����<�<�CS�D�7�(�Q�k)йW���MU�#�]�`gn�FD�[�5��đZ���7ۃ�p��Q������<�Q��ɴ��Z��%+m:��1>��v��~(2��c�ߔ�Ǿ�
��}���w��pR2�z����2ec;q�:�~tZB
_$o���W,e|�+��e!f�\���$*���;��0�Z��[`�}�(���X���tV��÷=���,��V���3`�,�w�����	�<p
ac�#m�u�y�yS������^��p����Fܚ�aD%T�m���a��%�.�d��#�ˡdANFjޑ����W���f�	/���Zo�t[b\��X��Q;}�3鴧�.c�o���*ޟ�;�9ycb����;<����F�����cW�S�繓�>�5T�Z��PD�f
�*�i��f�ٮ�f��rl�k$"��8P:'�Ե����F�_��on���x��_>�,��� d�pi���B��f��sU7�^4���~p�%�p0�8rs-AUy�*v��X����q�bP�$;L:����B�@��p(��f)ĶO dՁ<�����Tɟaq�>��J�V來��ן.�կ��wd�0�=�+�;�����?r��G����!�e��c	.t��`Zco�!@�y�d��#i����z�l<��T��r1prz����3��\(U3�B^<��悟��'�g��E�-��h[z��ƌ��Eyّ��c�7���C ��}b�g��>hԙ��{�Q$�.(���UB��~IӂD�rq����j�r_��Dt�/1��p�7���3	k��ݷ�`�l�t���{'���}Yn)`y���dew	�B�%/�`�p�ɞ����,��lM�a�&UQ-K[Ǡ@�*�-���|}9��Q��)�FU���8�럧U�Χq[b�˙U�䯉��Z�@���F��^�:c��.222���|�J>���ft_�&#�����*~�d�x�z���]T��'��OοG_���K6^i+��2�v��' &pg)���|!:���e�b%��X�'�|�1m�fu����Dh6������<�#,������ �~~���n���r�U8>�&,��7K� ���E�wY0򬪻�'��nL�TVNό�І�:�v`��8�P|����uQ�:��1r8�x���d޴�K]��+ۤ1tO��r�T'��F,��(61"�G��Lȫ���u֏8����`��T���@<2l�KS⹶]�N�(�`��e�?�H��O�C�e?�e�E螩�
Suk�ښ6 ��+�,����෨�}����o9 l�	.��f��3��_xWbĬ��{;K������5���I���TZ���7���\졼�+:
?����pE$�a��3S>�ʽ茥X}nY�Pt;�vx�C���G-~76.<�MVTQ��T*oI�ja@�v���Ͳ�羇��_���ie�Ћ�W/����St^��=>af�ޯ%��̙�E�b��ʮo�m'/���1S�!;��ty��m���b�X������&��2Q1罧)�U�n7������v;��{#bo��C0PCr3H��twz�@��Fb�^,z>�??�d���I�p� it��6�ǎ��#O��1S]������"Y �v�ͤ��cT����:p���7c�Hi�Vqד(H���a��cE�m��վ�*���M�����qoxӷ����{UEP*�nO�	,��BūI��0ʭ�!p��e��b�BSHG�'`J,6��O�������e���v�Lr�kmq��%�-4_`Y�,ع�A�QuODa�IW�OV�|�U�o��t��u6���8-4�)_j��3�=^��44�ۚ��ZgF�~S��T�~}* ����qc�=%$IV���(V2ֿ_Rh<}A!h�G�n�/k�v<e?��S�����^��^1�@���:�7X��Y(�ۮ��>���vD�`g��k ��ZHf�a�;�_���Dl9����;�B�î$���X.pٙc��2��P�MȪ6��6?�"��o��&|;Q�q-���F���$#�W%S�O��
y$��'`���\�?%O�z�"Q�<��ZZ���e�_�����F��j%�e%�������;����j�kQTٕ�0��`�
��ܰWlw����5�~���.Ʃ^�7�b��=~��l�`�������F���TЇM��c�b���P����lU� ���d�A�;8J|d��d�"k�d�7@CO�P�L�����2���)����)���
�BqI	�YR'�s.�ԇ�ņ$���.Z��۰�scF��ԝx�����w{i<1ۢ� �x���vHh�r|߯���K��������r�.<�pc_J�\s��Hձ`j�W�<�3S6�����X��/��[����Ds���}�X�nޥO4���7��v��p\7�4κ2L�ߴ	�u�v_���}��h�sFM����B)�S�q��;��%�jZx[g۰k��n9�c�[a6�2�R���X|@��2���`�����:�%8)����Po0���B;�j�5/����-�L���z��24�<v�e�	1Pp��,�P���Jq{�M�⿗p�hiE4^�6�#L��.t�y�\��Ò��}`�of���Aȱi�V}���#Mx����%j��6Րz�f~~)Y;�_�����ԮWO��~��#J03�\^*�=1]��C�n�)����>\F��˶G�ѥO!o��cJHU�O�=诬q{z��q�\����kU�q��E��$*>�*J)�,^�d�I���i�\�,�7�`ЄJ�Δ
`>O�8*Ө`y��Jfq��f6�"�{Ȃ	J�Fq}Z1d�]F-[��� Ul`K*��v�:/꼯Bnw�8��F���z����p��3�;e��!��*�}B\�B0�#��nԏ��D�V��'kk^����Q}��rMߪ��K��vLn���%3�*����-I�����-ǋ�ߝ�\�O33w��mˉ
�����_����=)n��?�l� �w~�0�Z�C^��z��Z.h����׽��B>�ʣY�:��U���!��/(.׾�d��D�z86Ex���1�|h�v�� %]�-���]~�&<�ICJ���י�,�.�v�\k#��d���n�Q3������v������=���3��Q����]ҸԞ3�.�k>�ez�;�.�l�)Iz�������	�QČ�DEM7��ظD��TT�3�2�����55�]��X2��n�g.���[۹x������8��P}�_>�z���� �NM�68'ѬX2�$2EN���{6��VhJW��O�W�(�ZC��Nx�$�D�����Cw~΍��]���d�]��uPHT�k1�n�Y7�&滧�z�`�e	���.��Vb�S
����$�h�6��5�^��:h񫆎i�vt����&��,s^�Kh�>�]Q��W����2���R�g�^�XǺK�Y��cZU�()���j�������Y�n�k�^#���3�����[!l��y^>3\�5�N��|��v���b#ʓ	�W1��2�����3�3oR#���HBɟ��_Ծ��nw����"`&���=֯o���U�`�I�G&i03���pֳ��`c.@�~ZxJ4��=�zk"����1I���}���TT���iw�c��	��wy<L����o�3���8w=$���i�����Oͻ<���X��vi72�j
�<��9�	��u�{b�x�GFSV��ap��������Fx#8iD;RgJ���adm͐�s�߮�(�N�`Q!ΰt�G�ɥ��+��ʊ^	��V��M��߉dӜ�m�:#�����3�5H�H�RD����ͼI�,�L.dW﬏���{�^z߁G���.F�J��G�y�ޤ��#�^�����o�ǒO<U���]��?`�����9�7B�4�V�0Zh_C��י��s�A;���	q
.(�E,Y�pӽ�ň�Ǚ=��QD��%UR>��y�fX7Rl��3q#
�1x+2)�]��U}��h��U���r?����}��.�a�T�Xӆ��ü	@/�C|)�+C�_�a�W=C��þZ�}�:<�O��\�]��*�5�mo���ֻv�Z���q�2Q���3*��x��wY��-������q���^Y
�=�R����A\�[N��N;`�%'�UɈ�b��.].-n��hE�ݵ�_�w�:��y(!s����N�n�H�c�1f=;���t�����"��=|h�����:���0.���9�̣��=�ܣ.<y�<���8�uzk^�M(DJ@�g��W�R�l�<���s������MD��shv�B��%�a���a������<L�*�T� ΅eہ]3ݲ`�'�IH�J�p�q���4^��E���`?����Ҋ����h���TՈ�!�aܿ����8��Y��f0�j[/6`���^�i9.&���h�����W��իD�g��s(�d�G�����q�lH:���iw{p-����mw˳�|7YJ<mKC�Ef	������������H�Rk����Θ87c����lZ�p2��Vkh@�)��9ln~Z�J�M&�j�d�*�~Ǖ;�7ŏD�<��ߺi83�Zz�-�\��xcf�܄(�xxmW�Dk�oa�D?f���jz�3��_@�fT�E��
�I���nBH�B�3�Vz��&����-{=f%)Cq��v6��8[W8
G������wJاl��ꢐ9�M�H��~�&1izU�Jyͯ�24\�F2��-���`��$�xq�[9�$ ��8�y=*��7������pU}�Q�G�����ȥ�����[w�;��R$��d�M8���������&y�x����=�\<NH�FbZ��/$$��:���>M�l��?�y�z�x(!
 �Nw�7�tH���5��oV1���H��W��kn�`鞝O��zD'�V6�z����+��oE���ҭ� l�r:Y��{Ck]��xd���~<M�;��]ӽg��|����Du�r�Y�v}��n��o20�gC���g�P�)t�MDv��yϿ�����(rf�	n
�<y���CR�Q}h����.4�U/��8�XU��8K˦$-h����b�j�n���.j$o{��qf�B�uJ�.��Hh6�k-z�=٩�TE%�L�D��� O�PP�<�����THt����^���=�4㑃73rZʢm3�� �d`�WJ��c���4�J��T�a��z$��֠G�����2�����ͥ�;yݵ�{�Z�
-:DU��=�]�qr�aC;�g��Jq#��7�E��C4��5}�9/Cۂ@e���Z'�����D���Z�%M��U���;�-)�םح���#�\��%��8�����pv5ɉ h�.e�s���hv<���clg��=��i�G#5�gUT���;Y�|=��c�:Ϯ���<���M�8r�����ɀ��ꢡ�Рߛ�ί�Qa��q�㐞�d�U�&����&*4}��)Ճ����iD-z/}���q4���"��PlX+2�Y��Z$��rlnѢ�)S���[?���Z�_��m>=LF`.�̿�c�:�B�:�D��BJ�0A@��X����	��n�=V���J1Y���ܲ��V������N@&]�_�\�@Q��b�5{\�WR�v���]�D��05I�v��E���W+���|��	��a�>�J�|�Tr^eE��qK~��4s�ͩ�����1��>L2�V�|V�9^b5�<lP��� A�Ex�K�'��u^��!�����xZ]� /���8ض�+-�~�=�?]o|���V&:%�u�Wn�����:����׉��do�3�i�e�܉���kn��k�_������!g�b`$��k<� O��`([5h�{����p^4���� ��9�����ه�e��kR�q��:a�E
���/gм����B�i�Q�3��#q�ߵ,��N|zK=�;|�A�]Zysn���4W��1	��E�f���et_�/֧�����+0�ibZu�)���C`���X:�a��*JpG�.����r�kdyҲG���+��}�B�&�E�ʦ�x�;�>�r�8��Y;^�$艞X^���/��F�yFP!����s�0p���P{GFaҺ�����Y��vD��ك\�W��gf�ڎ��ف���.�[E���������H�ML��D�JRI>O�6�D���P:;-|O�;)��S��BXS�th�Mi9V�i�M	nZ�"��#�cC��A&���ڶ�����0\B0G��a���x�ijZ{�g�x���8NX�W��o e5��|�:I�ď��������1���v\WL���l��[\.��Q���c�5�P�,���x��FQXX�5du��ЭܱeffF�1�d��f�$��'7b.\�eQ6:8���b\α���_%~=�
/�K��+���\�b�l髼Y��=H^�����{+�1=��S��d�aW����lmm_=����{�ʀ|4kɷe�K��"��@8g��Ͽ!�n��m�=.��lWHI�ޒ��Ղ���*�,�$CG
�#�g8x�Fn�5������Vh���D_"�?��a�3+)O�=�`�{6W��@�����!��xsg��A~,����3�B}�s���~���Y�h��n@�������	ʡIQ4.��q(��o�e^`䀬����������G����/۶���v�$U�2k���(*pIACx��B�"���*��I�Xg���Y�Ƭ��E�0��C��Z��a� YG�U n�x�S,|�˔���+�yʼ�f�W!ˡ�6�e����=H$J_��kS�ޣ�`���GC�A6�b�@���pTC��#[��Pꐻ�4��z\���	j �j\�}�#�!\xJ��W8V�T����P�c��,�z.@������wii#b r,��D_f	R\~�
|24�����q�m:1�������{�7���X���D��K~��U.6�w*��������2�0�gL�I���+Ս-��(��{8��Dei�9�Į̲���#��s:̛Z�vE�љ�R�����^�>��sO6���������V�!����A߮�
I�Q�����v�8���O'���#�>$�e��w�O�}��yÓ�c��	&��6U'�^�I�)�Vc�^������8�xrH��C��6���,���g�$�sX���'������	Z�<�fۅ���ڍ\[���9�A�WP�rn��]�Ũ������N��M3`\���da�����0�*Ng�`�#��f�|�Є��m
�,�E9����`d7m؋��Ż�vw��~1��3��׷/�Wth��������\ԡ|�>>����ۗ{Ξ�����P+eP:^02&��<Ƨe��tݱ�^�:���H��YU"m-�{2�L��,���N����C	�Qf0���D�� I_�Q� ��a3�������>َ;�����B"}Z�P��̢�K8�W ѷH4��h-m�X^��N=ȳ:۝Tb�\���+V�*����is�}h~A��5	���MP�F�UË��@��=��+iIq�`bh�����q�v�OS���R˺�FjaR��Z��\"9M
R܎}���h���;�cq7�����/�-ō�y����S�:af����^�x%��s=�J�>�=8�#��JWQY�	�ƧwG(��W��|J�zP]AwQl���wCM�}��uF�����H9DZ��:���^�?N��8��-}LX�w�Oq��zm?��u򦃦������:U���m���=�Q��:�}r�-�T��qz���~q~����Ti��7�rd��u�b�}�����O�s���̲��J�O���a\��e(���W��~���Q��}<��lbŽy^%(�0-&�����ZO^(�� �ˮ����m!��Q�����}����&�^��h�K���ɷ��d	���*N�l7�'_>rd��N��������2��䞧�tl�E"tH�а	�������YHb���ڔ�-T|��1<��g4��)>��M\(h�/_���^�,E���~_�H@���ux�ǿ���J5�v��V�N�_M��Q@ )y�@�0-���fg���������Lc��a����r�t�P& �8��HqDP
�K6!*�bo%|�i����9v
��V�)��R��<�k엙à+�&��c�bl[���M�f�N��2 sߞ��g�k�[�B��1��!e�3��ϴ�4���I��'����D]��%}?y�(�����k�ix<��.��ܫ��i�����	�>�;tf@��������R�VD�Ъ��ؓ|u%��G&6&���:���y^�������*�2����3`������tZ�a26�$�#R#<��'A"���IA�ȇ������<#2��2RY�P��Yk��`����� ��}پF����)p���>o����d����v���ᾁ�r��:u����Q*S���K��|��sϵ��R����WpO�����(>�0LjU������A���4
5���đ�YU
��=�	7x���j���x\�S��+�efQ�
���G��_��U�k�]S(k�:�M�q Tx�J�?���� ����;X�s�zEϣ%gb9��3�C��Xg���7\�q��3t駐C���B#@>OP>�j�_zw������b��f��H��[T�)d"����/�i2.��I��̈A��r||���!����ʕu�1,9�����,�,O3���L��m�i���C��FG�}Ͻ?>w* �&�����a.ZTq/�;/����{TV�hZ`>��8oH_y�ճ�`#��7h�^{��H:)�����kѤ���&���N��v�[z��.��(,i��j���d2T�חԋ˿6�Ϫ�Y���k���q0�i$�"���.�jsж�V��33�/}Չ��{Y,�ך���	�B�� �ih0�7[��� ����S�mzq&r���E\��pT�����M��<��ːab�#&;yb���F��.5��\��/�l���~��̲�%��FTw��?f9�M��@}m�b�!H�ܳ0���^	l�7q}�H'l	dfb:3�&�����_��XA�m�q��sux.C*�%Ψ��I5	�b�	DL����q���vXY0kb�P�I�ׇW����&�iT�E�L�I��([#��]��T:��ȋ���R��8�5�։���IiF��d�����6�������O��S�}�$�B܂�+�8S�]H��X�d�1]�d>�$P�VkTA3J�ul�F��	�v����b	?�`i!�l� -,$�9�5��/��"�@~�`�뻔X��+�ni٣h=�72R+�W	ŧ�Bx
�H�E@����a3����}:R�X-�D��3�dQ%�O�D"����΄�}��.P�VM�`-�����v���[;m\�'��ۋ$yLt"��P���\w��佣���Q$чc��f�6�w9-$�v/�����~�L�8P�o��
�yر����w�mv@�sZP�ZT�qzyp��D�{ܜ4q�@��滞a�{�±���nv<s�"�0v|���'�W�&�����~����a�`f����J��]�L��� �x�ڹ��6i��< plw�5ܣˠr��y�1�Y���r,9}z�1S�/��@e�����Wc�g�L���zx�>V75��� eV�M/ѡÍG��{�'[��b0j�1��8�.�|��JzV�~�N7��������/^�_ZP���R��BUOȮٹs��c~u묞��d̄Ι߮%^SUʐ�փ'�ْ�r������jXHE���7%ဘ/%5�������d��g�V*�
���떽Z��Էڐnc���D�y��68��i�!8�W�[�t�>&V�]DD�@e�3��fBj�F;7����*�i?�3����|j�	ByaO����'_g�u�Ƒ}���S���Pz`�D�[(�cg&���������ZZ��z���c��/�>O�1nW�r+�U0U%hJ��9�����F�ӣ�}�'�B���<N|x� �'�o���CKW��t�:�����	) �
c%�#kq�(�Ͻ�Ss-Ҵ᰹&Ρ2� e��%#����o�j���	M
DSCj�i����!T�[`����������m^[�D�í�O�ڦ�%sm:o<[��<�)[7fa��������������v75��! #e9��ye�R�[�����'H���������&I�rf�ll1A�]vÔ>���M��:8m�S��3�ʖ���<p?�,��Pѫ�V�Xn�T	�&/��V!��W,ʡ���W.��� �����ϔ�JT34@���
q��I�Y1��UD��μ�,i��SLU��H�a��b7�Tٔ�>�1Ge������J�I����qeӊ�Lm�)|	of�p�(�����$C�=�yUg��7֧��P��d�@`�&�8�^���D<�'�*(��f���`�t	��$�h���_/�"�m�I��=�&IK0؋&x��mf�"%2��uy�4�PNNN:]�>T�X�\#������$�i{�U�
�J����iO+^�������+kY�3��hq<�S���?������H�����H<#�L��ɘ1�����y+�Aa��Xl_�jB  �!<s#NA�4)�E��͎�@q�����T�~���2*a��+��sI|��a/��{Kc}ޥ)����"�)y*%;܎��]��N�����3QJ��U�6����#d2�������lc��F�s��@!�!yO��&w&������:����K�A�
�˵"�����HW2�Z��ۓ��E9�@�)�p(} [�T��?f�sR�Y!��H���3��G���ۋDh��tB��IVՇ�������،�=���l��̆
�72J5۵��-Tpd0��2$���s��%@%nԞ���n�z !�u��ۅ�/��ٱiB����0��&6+�Bl�路���P@F6ͧ/�M&ձ���L�q�@�2Y�Ͽ}B�NA$0ؠ��ȳ�w	�K .P�)̘w���:�4;���G��3 cj�a��7$$$n��j�y:�Kq5��˿,t��W���\я�Y���KrD�ذ��3�Z�Z?*B�fnp~)n>�H~&�O�D#.YoN��:���B J}D�
�,��l��]�`��k�Y
���� �)<�$�?�ݰ��
!�ޚ.}���5:{ku�

��g6�����&6}3���ϕ'�+S���ĳl�Ux�tcY�N�1y�tFű�΁�e�][O� �4��2�J����6ɧa�`��s�� ���0ߌ�;���i%�f}C�f�D�p�YҴ�P����ЛUTID�X�&�X�.�l`~ߨ
_^���1��~ҨO�R1���<L� "����N�*��4���-A�A��e���}Ʃ��K0�L\k{	Q��>e��Ao��O/��+�4��P9L��&"��/���<a�����5�'�ޗ1��[A��a��ah$��Q5Rʧ��O k���U�d�*������A�$���ۇ��#��Eq�5�F��fn+���%?iVE򶮙�/���_���)T���Z�"[�_��.)���!�)(Yܛ��9X���K�n}�ۨ^~X������-<��T�Y��Z��jO�8�"����E[R���9��b߸td�"|&��qs��;+��р����CA������,y����э�X�Ga���7T��H��XD��˻�[���t� ;}q��Q��?�h�&��f���ęi�qr�^��V֑j��~Qt��*�V�B��ߚ��/s={���һDݯ9�y�ƌlb�V�6������ȁ/;��u��JĦvf)�o�t^/�/G��J��L�a<PʇV�,����&�\-�����ḧ��0��������3�r�F	⸘��A	p'�BY@Tσy�X�r]�9$7�@2�XBS�N��&���+n��b��r?Lz���;Z�9��_<褒YG.ƈ����q%QD�С��h�kAQ����J�sW<����Z�O�Q����}u_��Q��zC�'�l�7P퍬���\��)�׵%��:�Z��u��)�E{5�D<_m�:��Tg���ۤ��rߚp�}\۰mM�{ɿ/�A���Kq�:|��P�����T��F=Ü� �����,?�)�˘���9���j/�R�z���ຢT��q8���<c):�Y��� Y�e.N$&�P۩an��d ��(z����i}����)�#�E�g��k'U�ݘhU�
��"AN�5�Z�g�̛p��+�w����8J �|_$:������Ts�]4+��巵X�57���!a
�F���ڌ_FҢZ�9���MAT/;o����F$������H+��8�h�c�a�vF����O�'T�Ws���;�$�T�ca����~%�A,��jii���fE��E�#�Io:m_�9�nX�Ob����V�����&�X���4��;�D�29��re�zX�X���3z�N�O;�������2�����!��L��W���Wz`�Ӊ$F���X9��S6?߷u,�ـ5��� ����~X̜OM:p?�t]��(��0��}?V��U�N2�$��Q���Y�Ͽ׊�{�nnrVj���kv��!���ʺ�l���#���:lk1Y����F7%	$�F����0�r�����>5���İ	�7\E^ȩ��Ek�n�u^�\nNT��h[�~�⓰p�򎧭��jb��ފr&�x���������d�!TM�s���؂�-�z�4m����.,�$�EB�k�����8;���q�����Đ��b�����I�Z�|��IG��.$cD".����e|�{"��N���[E�1��ZU��dj��x��v��aM`�F$~�#�����l�}7���#�G贅yf���7}6���J��.��V��|�!�U�m�wᣘ��m����Py�h�`�MCI>Ռ��� ����3H���gڹݒc� �T�1��k�]��X�t����T�>�4��P��g�ָwiwI��L������;����Zx�S�ϼS)���ϗHS��!#1G�\�{�t�܁��]{g'r(���R	x�NE�����	��sYe��+�bbc9:�qe*�����%��\l� �����Ե�ȳ�Pś.%~^<sש�`�������n�S��0���RU��z]�J���]�̋pg)ʌ���V.Z�<�a��>"�lC3��j���/B�B����B�����ks��t�1�ԯ
��w��(�S
��"��Ŏ�k1��D}�0 +l�C[��-��f�$K����/!�-�#�y�19�
D%l�c�CG�k7u�4҇��"?���`{/6wM�i<.̼�h��G^eK��"��a�I���7����|{$
5�{Y�g�l��,��!�cbCi�P,��(����;�����5W�lEG��E�/�/�y3���ˮ�<?233Y#ĦC�]LQ�d�-2o>Ѯ�D�&Zr̯�q?�	6����^0��C�2,ϯ�+6h�</�^���T��$�F`������?�@�3tp�|�yR�\��I�4���b�-�s��bz�Q{7��9[K�-�N�O윩}p�Tm�(��g����I��J��ۤ�ƟW�bZd$�4�,|'��[�k[���&ҋ$v�w7��"'�n}~�r����3+QG���kT�y��4���C�p�y�JvɛZ�l�Ĥ���a+OE�v~)WD��J�^c�]��$�����M��X�D��dv޽��~�z�z�5v�4_��Ũ�0#K#R���^�������[�n�]VmQx�g1�0?E��ߪ�V�o����O���'N`[T�0����h���m���$ä�G�����x�I����u��آcE���;}{$�p�Ob��k4%b=��	�	����=BM�]�
�}��ᬡ���h�J�>@��
�XVjQ����B�m�����~ۯy#,��Չ�r�,��>lb�{�y�������6}[�j���������w����C���y=�x�⌱Z�pWXG���4��e��8Z�u<'r0r�AZ	��"����`ݎ ?G�{6��O��8�J�����%��*�������_c@g�Nr͹q� ʧ �ex�Ɩu��	95��������H�)!���J�X�G�܉9`��
181QB+2��1�r���Q�_����~-�	������G\�@a���1�WWX!d ��w枑�`?�eS
p�6I��ߒ��[���&�,����1h~��˓ �X���]~�F��g�ކȄ���X:p�a}�P�_e�0k����F���9|��"G��� ����?�ч���Gڤ>6M�����B�s����K8i3�\BB��Ĺ�4#bX%��u�.G�?J���"�7D%��<A�j��jڦ~~�'�eq��<��C��ܮS�K�C����%�ూ�� ��o��r5���"�g�mN,�[�{��λ{�{i�)&�-ٙ�\���Yxa%1h���q1V��i�U;)�����Z��\)�6���F��I��1��v6[b��L|"�B�'�։ĕ<�a�tVHl/)����6�}�L�
�540������/Z0�Z�_Ilny��&0�O|�y	M7^���{��{�Ǿ\�r�ߕ�	�w�un"EP[h�ϋ���_P���#�ZA����^Gk���<~Td���?��ˡ�=n���)2G.m���N'S� �;�!"�&���+�r�cz�#�㒔~�-� A% -��PMX@1�0�R�h�̸kG�w"�_�Y�Z!�8���~�#��Hf[����8�s��O��%[sI1ԌEI�E|�r���e7��*�)9�l|
���V�_"�d���׭�}䎜o��"���'�O_�eP��A.��B�8��E�I�J�*��u�^�ߝ�`M/��c��`�Qh�Q��^D�=������צ�V�FI$�6��V]3��X�#�����b]�n�̝��K@��+5��t���9^dHg��̎�N��ʜn����o�5�g�~p�B�ˇ�'!~"���y�jWԭ�hQ�����T�8Ɲ��B����Fj���jw����l�Lȍ�DF>Ϡ6��8�]���>��\ç��䦟9\-�~9Q��ۘ>L7�IČ	�)������RH�C[�f̨�c�-+������1M"-
�&o�ɞWe�wsS��ԗU�q�y��SCC��C�M�23���b�2Œ��h~Jla0x#��q��X�1�e��j��4P�ĕ�.��%�7#"F!0���J�"x+�R��_���a�v�O�
�r#@��@)�̩��k��	����� ��Vl��I{B+ǢvE�j;5R�DlY٘�U4&4<���.��+=��F>[맾�ج�� #)#���5$���fG�$�8�FTw&<<�+���\߸6{ה	�0�*��&����Y���+a�b�G�\��XT�a=���a� ��rhL��9��ĸ����d,5b!�v��q��)��L��KՔ�7f&�qh4.�8z�].%*���'l�]��}�{�A�z�*:gv-#`Q�����l�zW�݋�I��z�iq���� Pݴ� 8�_���ޢq(��}�7
k.�P�p���䌩�Q�F_��2�)� �����R4�����@8'��F#�q�Baj�S�s<�s�wYy���nGt�N��S��L�6Lj�{�ϑ5*ɓ}	�̜L�뱒�7�E��&��:�r���uXo�=nj,u����RFH}c�XG��$>>2|yf�����=�|�/�1��e=�YxK͊y�D���m�����L�lm��n��0���vM�nl'۶m�ӱm۶m�c۸c۶��~�Z�>�����q��s^Ń��m�R�}J��JZR�s�`��42k��<oΚxC�6!Ieq�g����wf]�д�6
FXV�.�Z�R �uf1���g�+�7��9�J�=�?��:,�����V��,z�8����F>.k��	c��>�4*�l.���A��Nt��N���3�;��GD�C�������vmWˋݙ���ͨ35�,m�����r{��#������Nea�<�&u
L,N�w,jjK)Pǯ�.U�3E|<3C�D<�@��M��"lM��g���a�	��i��*+5Gd*�w%T� l�6����"e�7�������J2����5|���6�a�*��Gp�2ٚ�,�j�ٓ�L5��q�W���9����or<ݧ�����H�-,Iw�3yN�j��C�S0�W�1*o'O� Lq<�j�$T��P�kQj�S|lS���ېCp�7�u!��7�t�����3��C����Z��	&�}V��Ǝ�����Θ�#������&�й{Κ��W�m^�����U5��t��;�7ΝΛ�מ�;#@���-u�4�q.y�:��r�
��1�?N_q���:P�yT��zZ���R����N��Ē�Mg׿p�h��B�^�.�J]p��U�~2����.]�<���O�G:b�}z�T��:��#�A�c�O�Y��"��*W,V�'v@CW��}���Vր�<Kr�tq(eP��,
s���SJ�p�ɤ�����32	H����u��0/��j.��@�O<}�K-B��B'��
�p��}n�x�_sý0����#<s���i�S0A�)y�f�j����B/y��a�
t��ic;M �PY��Lˎյln�+k��~���\1��P	�%pBR֥�U�4�����L��{��Y3v=ܴ��m�^=�ޫb|�s�U��KR�^��C~)	2m�kbm�β�Ґ%[Ó��!0��ǵR3��(a^�h[��B��C]|�IH�ЈU2j����B֨i%��Y�������X�ó%d;@�9A4�A�\K<���͊����q���$�+�ԥ:�VD��l�6�����7���m��,~�D#=�俣.���9�����q�7=7�ߗN��2�B٤�-,N*{>g=���}⤤$Zz��ᴞ��y�#������;����a\m8�ή�����\p�� Q�P�ԗ���󶭃��N��	8��+��v����=x#SS�Jr�&�O@��⼇�F�i�p��-O�f�N\���#)�XC�V��Hut�WB����/g0'��d0!��ب/�h�?e��I�R�:�!��+ȁ����C�.���Y:Mx�6��襏��u�hx�o>����(�pE<�45we"R�z���O��sE�gG�E�K8���3���.D(��I2H�Dg��!�(�8��u����	S"����P@$� ������>ׅ��D�ӌ��I�L	 %�YUE�D~��c���,�i"��q@�>��Y;��X9�T�
dU�H*I}):_�H���-�A~���ÕG��8�	-}�
^���U���	����=��m�&Α·+a�Dayu�����%+A�A��|��5��(����q $�a��i��v R��KO��?�~�e��m���ql�&�r���!� ��Z��;8$�3�a�h�В��`���^$����m �Gx>}&W��$L_"���O��������v�H��Z>���o1w�$l*L6�mӶԢHI��Xy�0!��U�BE��{h};�� �pe�lˊ. ^�h�G�fU1�~��wLUnB�i���+���3�<	�8m�l^��Ve��>(�|}�R�J����K�פGv�(R��P!)��h�5ђz$sZ���l�xc_��qwPU��x�^GƁ@��
oM	 �W�_5�B�g���F�1�N&�6D9ݏ3����,��t`R|Q�)[��h)���&��`���1�����`��Rm�#��PU�m7��H����1E������[Ȗ6<&2��"�g��I=�O�Z�x����H�}���|b'�;�ת/�]֋t�0iй�w�/ׇ)��t?ƬТ��nO�v��iC��f �ѓlJ�m��]���&ҢE5�s�1l��9ӫ��o�_���G}������R��K�9�3o�#�V��"�i$uI�_�4��E(����gqM4z�a{�Q�"U�*���c��}ģMa�#n�E��J����=y��qF�º:�����q���D�� �&v6����?RT�PD��F��B�w�
��,�������ٕ4�����	�扃���P�'�$i�ၽ��C�y�@{G!͢
�A���O�5�H��^�e!t�/��`��\f�*턜Ų���夡�������p�cC��u�����<e������>æ��s�����ieE�Ε���\�c*�����/�k�L������|��/�6s7R@r(�j\������c���k��S%��(>�7��-�G@2�ǅ2��Z��/,:Y��� ����u�������OK���u�Ia�>2�69y�kR��t�z���v���_�2M_���>��7r�렯��Gmj?�[�����	�y�M`@_��H�}��BK:�AsU��)H��
a��N�G�}I�	�}��-Ox�� yW|��\=A���/R�2��>��w��d�f�p��.�_ZY�����|r�F�=z/���i���0i	��3�&�ת+�%<Qg�ԭy}�4iW�"�\b�x]�nϢ3�.^�����r�5��f����'\��3��b�� qVr�K07nF��p�g�H!v)�ee�v=�kp 4pdP��81�F������F��(��
s���Թ��\=�%����ʙہK�4�UȄd˥ES�U�{�
�A��	ۺ���*+]�s.M��E)�p�ZڴW��F�G�(�Ec������'��OT]�3Jy3�>6э�R5��@��6�t�꛺��5�qj{���w'�Q*c��f�Rű���A4)�qLU@if��Ⱥ��]����h�574���!��!�i���L3L�'ٷ��sLݍ�����2����������i!�"���@̎����~OӨ���|}���q\7@	Ѡ��~~pz?Bm�ڙM,�6��AA�x����j�/�J�&�ok|�����T�y��qG�9�3��Z�F��?��A�"�vQ�rp�ĺ�@A�% ��t��Iy=��z��av���MZlҺ�	!�/O+��&|S�ש)b��&�7� �=�m�6st�6m̨KJ�$K.2g�*(Y�aGy�g�
��|���6�-��;���\��?�� �ǲsM#+�
!g0>��QR������b(�Vu�}� �^��W$�����O����a=�#.!N�
T�z�+�i���K�����P�����{Ï��	B�S�%)uIZ����g٨��yi3io�:��K;�:[�6˘n���E��h���j��w���d���:����)ˠ�o�^��X70�v��墕\,>�tM6gs��9̎�1���҂���Y],� p��/u� �H�ay�-�8��Q�y���� 1�1��F
ӡ%؊JS�y��IB|�:|`J��B	D>fhWC����%�|�N��+�K��3@k��+v���s*d:p't�)��#))�5s�z��FV!��h�j��c�����q�W��͝�gK3股3]s�̤Y���Q�f'H�,v	�b���0��nԧۖݴש0����aYU��*&����A���$7�Y�USN{��i��֨�a`�(���d4������am���׎�A��vc��oH��3��� ȸ�NᓲT�� ��S��T?�nM�F�O��Ѐ�WӤi�ջ��u�z����uqui�=�n5�	�m-��V@�M[��S �V{Z�C��	�����y�^%&��ׂ>-*�mK�`\	M�l@��.9�_Qٺǳ�A����*�j�����~� df�����/5'k� H�d��or���dz6�x���a��q���!
_�>FO�p�����Hc:�eۂb��_��)k�,c�:<��fiz�L,��>M�����!�Q�,@a��Kf˂1���8���h��m৫�+���o��z�gz��I�?)�{�����&��W�8)�n��0�Љ�*��\�R��[ �޲w������(�Sh��\ӻ��Y�qw�B���"�Űb $/�����w�K|�� �z߇;Ng�a����g�&q�����"Pikkٹ��xd�pv�4'�ޑm�o|�����U����گ:��:O\�R�����Gj��ڨ���P�'���_�F���T��Ѫ�!��0���9.d�&���TT�fI��z?�^��L�^�G �j���6{ӈ[�!I��E��l=�1v��b6p7N67'1��xi��kC.:�+�B1qt�k]�����Ч �g���/�,w"�:���`����.��C����uUL8ܥ�������3n�U��k�K��7|���d,��;ф���+�'����c�#3Er 1�nFp��X3H»m���o�	x<��w�^m5�H���Q��sE��q		(L����9�-��v�?M���#����*b��8 ��U]E�QZT��K"������:�H1�}U�[:>��𵍶Ǜ�v��u��7�3P�)h/^]�e���.�f��fH�U�u�0�Bϡ�hD|q�uu�I��G��ڰS���Q�k�J��G\}KG`a���u`���*N/Y���_�Y-��PqLԋ�{�����<녩jH�#I\�0D�l�(�*=�*�<���~���B��i�Ұ��B�����l���B�m�Umi�c��,	x�9D[�=��Pm�=�u��g.�H�'j�B!w�6��r�9i��Wb�w�H�=�h����;ԋ����EH_@h��}�I3*l��'�,6�W��4Q�"�E1���;b��B�����;̝l��B�T(=&�7�}eB�?S��)'9g�}&�-O��� AG��+�r� x6�O`}=�mϓ�����om�'s�|���cpD�:e�����[�_¼dD���Z������ iak\@>�W��&)*2�Zq	K0�vR=�!���F����s�ޱa��-/8hؚS��|��g������)]�?�����,	)�z�ky�	1C}�/��:@ج���?���-�2)	�r�^3��G�ZR%��j0�3J.�������b������KЇ��$�xe�:�G�x���G��m�O+�Ps���% a(SS�rjI"��t�UH<&P���v�ҹg.'��Yu��U��f���h�"�jU5�]��d�#�hن��IT�޾ D�~��^1�OA��yN|a�+��>(6 �q{ݒ&�#��5"_��z� g�G��p�>��\���z���j��ȰҞ�`�*�:xyP��ԫ�ɛ�E�d�5�v����h��D��M���o���%a��7f��Ȝu�>�/�+��i�M������J��i�8�~�ξ�%�v�Q�?�H�s�)�̱Z�Ri�l��U;%:"��ē���
�ȋ%�Ud�l�㡈��#D��Y������aQԋ:<#��L[c^
eV�X�k���l���j���z�}����p�Ԥr}��q��Pw1�:z���V�_�;v�l+���G����7^;�th|F�4 D�?�E���DeJ������-�g�%��죅����<�����KA>�X�����	��qT�./��	�$I���ց��a��HCk	��%N|nz#�1RԹ�!j���;v�_�:��6E�F
8tOh�>��w����<c���)��`prj���}���;M� �9C��p�t("|��0�J�Kog�i�.m�߅"k�`JAٝ���"6�(�r1��{c���$\
-ƭg��yq�sNx@�tw#<�F����uL�}��r�ˌ�)��O}�	xEC^��;f�� $�(�4}��Y
Q����hX7c���<�̇�W��@�����&��t�-4�D�	��$?3�Z���O�e�a��ժG��trr�Q��j
b��69�?O����`TJ� ��7�OZ��H�
�r�Ld�M=i.�nhQ�'�	w\Tr�ԈDv��9�G�^e�#�F����1����ӿΖ}`״��'?���s�"�=�?[�B��b:�	��s��	�ک�����碘��Y)ޮm��XG�i
��x{Or�K_�����a�;f�7:6���s?��L��K��*��X#G
���q���+��Jc�[ڸ��Y'���5L����A�C�*)KW-\7G,��$x��kΊ=�<����Y�������td��,u��p |����8�I �9_�����e�U��pwS0����b��z5� l��
�/�f�ab�F�lN������U�.��n�_+�d^���d�����̌�(%×e)z����I��O�������Kq$��r~
:��F��S��xl~csg$����Jd�#fv~����;�2����ڝp{��A0E��9`m�)_[�:�4��z�k��-8���j�gf;\���$c�{%m����e\��o��V�)�z2F����oS椹�A�ɉtc�t|ӡJ�0�1�)�%��P] v���eݔ�������'u�J�9c����Bf�ͯw���������Rr������I�8���Eҕ��Av%�5P�n�eA4��u�+����C<�
-eJ�A^��_?��[���C|�R��F/��s�W���ߣ�d�U���|9_[�}7�;+�Y��>��`����r�Z�l~��1C��N���p3̼m��oۣ�}l>�K��<C-��!�kq�$��<���0��^ۼ0-"ϻH�&R܃	���řvƤ�"'NW��$�xy�߉��i�{�/J��"#�׫��#i���>C �[k���JrJo�@�ܡ����i��}G�
�}�C0� �kI���2���鄏��F�И/WI�U�����IxEJ��`/���/Hgh��"�׵Z�BYi�Mw����9�N���MV��:�U��H'�6��6e��1��7�A�߇��ʼ�w�R����KT@:E(
�<�$.FG����H�m�`�eR�p��U�	c7!Xߗ4_m�1��cJ��C��[c�W�,n#X2+��'[\�qM4*���p����9������Iݵ�������mp> ���;p��>�����d{8;��ݮ__�f3���R�����=�v�>:3�3p�L�!�$J;�SU[�Hn+F��������^ַsKJf(Wy�<���|�������A�鼞���+���SquH��.�\<q�s/�iN�f�l XT�(�
2fHʔ��s-��5�wh��lnd�z��S6�������(�;�:'>����� ׳Y�;l�����$mV3i�H1��.E9�$KRf)t�uぷ8Y�S*�H��w�azPp؜j?�Q�|#rj��]ħ,�7Y�G��K���'���9�uד	R4FV����������l�s�U�Q�l�y����Pa��1)z��B;ڋBp��I=w��Y�ȉ�G!��o�1 ��u�q���s��5��z�_��Ԁcb*h�eq
=�4(�v\<yv=q�;T{T�1�4�$ś����AsD��#M�fdc+[(��L;��@E�?c�ŕ2���!�D��ײbf�*�B��PE!�!.��ˏ�)V!A$ a�����eQ�R4_� <��/q:v�W�\��7�x`f�V�۸L��f�oƘs��M�
�Y���aٽq��ş��w����#���йT�'�#.\W�3J\	b���K�v�PYj���x%�zEAl{��|�4a�Dy�ݳ3./��އO��j�ϻ�x4h�1ލ��E�.�B�4� �p�El�&z< 爠���h@!�(2�6���5-p5|O�N�e�!�7k[��a����/��G�o&���V�ёyeiGo��4�[��<ݣ�})|�G����,U���36�1֨�i��W�ܴ��j�X\�q���z@��=��
E��;��m��_^���L���I�I��;�fW��A�(��v�s��=��'�Ov���7L+}�̓����
S'��Y���3�*;��l�p�5>]�9r�*M��/�s3&qBQ�,Pe��_�Z�'mT�6���{y_~�?�q�)^3��"�z�B4���5��Kz_|_��>�{�.~�/����{n���b	x�U�,-#�r��c.��4�(N�X��$��IQ���<�#D)#=��g4��W�"���)�]�		/~W��bP�/Ӹ�S�HD 6�~�(^y�i�"$#��^�s���u.>�WЃD�i����
�
^3>��J�����tv��O�K�[AC��%�����%��Sx�%��x@�q%�\��;��~i��*m^67�-��3+>{�@���l(� �i���R�b����7À�^( b�섪���|�:{�L�G��t�+&n"��mb����ҷO:>j����Ɨ�r�,�͉RL��(->�g腯�^�N������4�G�ܶ��̦��x�z��9�תU�P��Mͤ0ʠB 1��(�PcƼ=[N4t<�=5>&qXA�Q	Jy�I:��ʚ?��S䠡2���~�}ة�8��=���4Ί kZZ'[jn�i/:�fp��2{��׷�A���ᙇ[����Ɖ��N�k0������c##��E[���R&��m�|���#nڲ�}2U�m<����&pI���fL��)�l[�]|J�Xpi��^G�h�n�3>�%Q����c±̡�"�xK�C�z�>�9+��W�C�	6�L�Hr���r����RS���u٭�1��]s��'>���8�dp3�����z?rv�6��r�.^kR:;�./S�n����mϕ�Y�w=C�v����&�<Hddf�7kY�ܠ:��^8�xDh6�"׵�/��T��j͸z�Q�-@�͞��U�k��y�^ɇ��ze�,S�(l|����ˇ�|��R�x�r�0(�>_�Qd��9��}P��K�� Y|CX?z\\E}����������Q�h�'M�ں��C_w���&����E��6KgED@����lny]��C��e�����x����0�{���`~���c�`��WK���94l�j9}���
�/��0H�g�������@��\�X`��S,-sQ�r@ㄟ2�Fχ�F~"�$���#
����F��{�:0�W��҄����(
��E_��[���@�n]�,I�8�촅�,�x����
S�_R�����CP�m��c�<*�	b�q7���F�\�*D�������wJ�+�h�6��W�ԉnU����}68��bg�$����Xߤ�'��+i�6qy]�G=&��K�y42O�}9%BNAQ�8�24��-S5.�;9%�c�O�0Ɔ9�D;BG�4;ԉ]��b �j�z��I��M��4O0:��&*_9��IS�I��(
�JX����̩p��W�`!'>�jb!��ղl��nS��>�4^�u9�c	�N��ޯ�a�U�?��@�P��$��R�1�����)]/o������{�y�?C3�$�� �=Q�\�J�hҤ+��:I�2)�T�5:]�������W�./��,��� �4�ȨѦ�����I����&`慒/f�X	���ĖE�JNy3o��o8z���`𒝻0�167�a��Û�����<�1�;G9��}.:�2I��T�-nm�{a�g�|<��g����V�ӂ0s��3Z'X	Wᖖ�Y��O�Y�`	�Tq�e�P�g	RR(з
ł*�nZF.oB�$�iT�{�]y'S/��F�i�pĺ�[��*3b�<(� �R��y[��lna�;���ə���kJYY���K����~�Ι����_���"=����W7��Mc&��C��Y~v[���L|NO�꺺�A���&&X�tŸ3����	���H��Jh�`B
:�4ڬ�u͒v�2�U	�E��m'a����֬���{`L5�WG�;� �`����BH0B`����~|�j�h���P�:��q�����s3�cq�Y�1�S�\��|�+;q��<YU`�[gL)ǻ'SD����.%00]S�>e֜����ɧ�H���	��B����|
�(���ja�:�E��.Ⅵ�ў҇X�@ ������|v�(�"7R�/@��ʠ�0��w dv���!D��OC��/D�i�L�	)�1
���ú抅�eb�R�N1���94�t�R�z%=/�����ԗ9�9��#`�@�V�8�����%l�YW��T������BO�3bIC��TN�������Ǜ�U^r�(g�J��	₥��gd����YӜÛ����Mf3���9��%|�A��Q���D�kGx�^�>a�������W�Z��t���>�.���lJf�����6�<�va�0����QXΞ0|�O��N��^ɒ��q�=K9�&���+$���s���h#8��L���oЭmF��=���������?ܞ��<������/��7:)��b͢�E��]�S��"6�X���]cO���;��Ϧ���̴R��E3(���L���Y�?���V�[C��N,.�	C��ދ�>?#	#�}x��d�(1��-A�8�p���p?:R{��y��Ƞȉ?\�t����9�������O{�,z9��ؒ���H���Zdg�ʤ{A�p���e�O�}�8��rIU��_���Z{�����Uw��/J����O��z���t���M�'B{xx@#�a͒���̖3ƃ8X���$� ¹�+�����EB��m�.��i�������r�o�߶%�� � G��0Zr+�p� �+HV�yٟ��{R���*/�7.=�5����jJ|wÖ>ōP�#��:��i"��������Pc"�#A�M-�YĢ>���������M���fm_B)
8����oH=X�g�ۏ�Y>����<1䦍���~(�ˆ�������<����%F#�8�"#��xǓ ��>Έ\��ؙ����E�yQI�KlMX��7R*�����n<[��!���y�q�(�y�%���wa.̊Y��ђ�/�fU�mТ}y!#%�B6ck�y���#|I\cT2a�3��"$�K�a�T�dP�,+�f���A�N�����^��go��c���{^�	�Sk�i&ߣ�III�

����-���Z�X/'�ݾ9��S���fӛ�A�|C '39'<;>[�:��\.�h@S�A�����%Rҿ�������4li��V��J��ub�����K������0����C��������a-�PA@X��j�O`Vy��w!f�G�Li��O�)n[��+zW�.�1�!3Vi����x
6�N�yCG�,s���M�e��L�B.������pE��7�d�?i�,��Q����q�&�7N�J��j�}��%Y�l>�uM%�,�3������1���!�{��e���s��Q�#���avk��܀���7!o�^ǂx?�Ј�]1~��i����.5�x#n�����Cd�Xc�h�M��j�]��A�z3�M���)���Qࡱ�s0-| ܛ�<�>�h|�H���X��0���թ��"K����+�>M'�.U��r�.�� ����S��.ܸF
���f�Z�J:�}��t�z4vm�����	�9?��|�	�
�v������ ��H �մ�Z��Yi�yr�v��Ð�[W��D'�OPHO�l>��rp�š#7���i7|H��Q����FEAK����BZ򵘿��~�1̠�����'j�D��MqT���q_T�@�[��{f����F�B������[��3UNr8ϓ�f��+/l���e��`�:�%	y��5n@�{U]���=��������
���{N��MU����g�gZ�9�1�=B�W�at�-��1X��`�z�*n��|5j}S�2���Rā�I20��rcK;�it����5���t��ġ�h�|��Yޘ2�:�*�$��ڤ��1�����Mf
L��f�L�����n�I���`��W��2y��C�1�HyL\ߛ��o��x����2嚻�#W�ԇ����>X��Λy��U��!�խ�"��N������X��\6%CO��2�.[�u;M���P��9Usm������n�k����>��J����سV$���Ca}��?Q�^i����}.�Ʊ�����3�Q����P�>f�,{ٔ�jL���{�覥�R[#a ʜq8t������Ϻ �x����3RT�	��Y9���M�����T���-ڪ0��m���6�r��Tsv� �su�n��/��f�X|37�,��؇۠����]�P5�W]�a74��-�q�֩:�Fj��䂐��}}Z";�jI�RbR��ҳ�u���Z������<�~nY��m"tiii:�l]C���
�����.7���>�[�&!�E�nw�I;)�.���g��[�,H9����{�L�:��������О�n�V4d�9��:��(~M�s9���Ab���T��z:$*)�G���v;�S#W���G��D�����_7�L���A���$�+����:t.W�8G��A쓙��IUޣ�����I��,�!Z �N�Pl�V�"�����p��Ʒ�g���<X��_q�G����Rc������v{�O��R?�N��2:̇�d̀��v�2���-^L�n�v� �ej��!���ˤFd;H �\�+���w�߁��x����"�@�r�X��Q�j��4V���y�Z�b	�\�׽ <�S��:��=�om���z��^t!�R^�9�+��� �����&����ܯ8r"@���'��K�ۑ��Yh��#�� C�\��θ�k�x�(
u^����
�w���vǣ����v�U�`��7~4���z�������a�w	e�t��
��խ��ݖzx�s�a�,w/������M�;] e�+$ ��_�圢'�զf�)�!:`�s�n,H�*<z��>d�5RQ�����-@�F��D��w����Ư���F�s���q�jٮ����n*ϳ[�h��HD0�������z�)�y��[!q�X�UoYS����C�^��<̹��������u�uy�r�j�Z%UX{c}��}�����'.g�N5U�m�mrd��l&�(!����.���c���!�j�$�|��ܵe|2'}�7v
o��2C�GT*����c>�,��0&�䬉�HUr�t�X9ֹA���z����L=#_�S��}���~����OɆ������(�X����$+����H�B�z9r�p9"���'B�q�j�X�i�\���G'^_BK�£��p�_�%P��{��9�[�A�1��[Ǘ�(;Hz�p��z0&ר3v�=�ug��#P	+��L��1�⮽W�;�V1�8����L鏑l!!���8-&���(��I0V,n'#Bw^4�b�4����:���łmMX7h��$/��QPH���zAE:r�;jol�����f�)�*��W��N����X�Y����>����	,�z�*|c��r?���>�\�	��� sJ �H*�'ʌ��+,������Y��瘚�vW��G�t	��`Á���9�x�ך��֎�[m�t�t#�8����κD;�x��򪪌��T�C��-B� �鯫�� p�Y�u|��y)¿^���D��E#[y٪�B�Y����{&��Ie
w�"��z��
���w��ß//�/�3bܞ���	҅<��R�O�2T�o�f�NWAV+�18��I�W������*f��5�t؃j��rL��i�Z�H�4�[%�g &�y&~�����(���!�^�������> 0�㐐�824�!�o��
�[��=�fO��YV]o�o�=�0�8K*q�������l�2e�~ye�|���8n��_��u߇.�,T�e�����w�7�)���~ �~�ZI��p�b��}�pZ`�q�'��m�8��,���I�3\�2V�|�Zǃc9[�j�t�q�z�[I�HS�<���
�v_��
��L��! �ý/�n0^�	Q���{e$��V�ׅZ�����O1�.Q����!*�'UUUw}�LՉ�����:�}��^�@�	o�#_�(�2]ƺ˕h�-�ʊ#������&�x6O�-�?�Gr G�=9.�g���o}I�$b�k8��=$��.���ٱ3]��Nѱ��ߒ�2��dmC ��T���@	.߱��>x�w^ƹ�E����$#�X�o�@����5�W`J+8h�x�S*1S*�?G�Ֆ���%R��,L��xf�tǧ2Ra'3�B��̧1D=+砸teE�1�}\��C�,w���`'�[��__w7��V7�[ ��{�q�P�PӶN ��Qq��Dᅖ�$�Nإ	��զʘĘ?�������֡�4iY��?��@q����h�r�gd�2)e6�d̙3�����������YMh��f��b��I����M"��&EF_w������ �Z$����h�&7��W��F��5��.U�E���m�v����}��G��!�8�������k��o#/�T��>;7�<媛k�����-[�Pĺ����y�q���B�ч!�������?�㿂���04t��ڤ�H�o
��6�!��񊠉㷤A�F�E���c;�ƔD|�\5*�Բn��v���� H��#�k[��0��`�$|��AuX���A�G{�=,�����)�/�w ���l���,[�����؎|3��_��y�:Zbs:_$��z���z�����=J�4f����������Y@؝/���1���®J)�'q�9��-VR'm"�)Z�#��u�p�[���ɿ~A\�8B�����Kc�l���>���$�\_.A��'9x}�p��Y-L�����H��t���o�����,�@n
��'���&��V���%7��p���m���r
o�%�x��D��E�u�K(a���ٳ���B�f�3)h^q�؍�����'��?��֗��}\}r�Y ���[.X�/$z�/d�+�8�ĳ��h�g9�m�3?���*�Ҥ���2�90!����%�{֜HVK�/\��3gdֶ�8�F��_��7�yZ~gI�9��Nu�ߊ~N�ȋ��m^ԁ��h<tܾTX*����B�Z���;Vi��k�*��5QPH��򳥨M���:'����u+܅k�1�w�� 1"Z#������\�Ў�j�H���o�*\��B\�9�q�}��b)����$e�dRވ���V{T~��7�g<�#y��C>(�ܱv��3�f�(I����nS1
�I��G.�vV��k�_M(P;ZX$�햕�b;z�"����Q�+���=�[\V'`S�� ���I��`N���)����ؠ�R��������+t�#<���W��O����2��f�'�uo4ڍ􉣚��A���	=B$��Z���j��Dttt����.�$H����f�]h;w��}n�JPvޣV�/��ɠ�A�c���˘0���F�5�$ц�J@��d�ƫ�={
|b�Iǝ=Sfyޑ���B��Uv^^>�s9[&!Y�wl�B��?0=1�o����Vϳ�PyӦuDS�}���v����.Aє���,д)�&���t�,&��l��N*���*c4ns��Ń�pZl^)]־��
�fA�(�m�g~�Z3��4ܯ�p���e��ȵ:/��w����ȥ�bfh8�����ڭ��Ve[����v�y�"�z�!:@�G/Iz����^D�EU�?�Lɀ­��W��*�P�>Շ�C��S2і&��Gg�\)9>�[�bN:(Xf�	"�L�+�liΞIH�Gi<[�ǖ�o��I�8���3IIqQ���3h_$�r5����r�o�����og��V~qx-�0��N�V]�f����J����(f巅��.76oS,���sX��?0�QR�E-VΙ�	L�5�i��j��u[*��`�{�2���q<�u�ޙj��>
\�A��� T!R0����6@�k�aJp�;��f�-18��6e�-��	���(Q_��X7���ӣ��l����,�6��A���ɹ��<�e�>��O��I��Amo�p�Jxt_
����y��Z�G��C�9��m�MҠIc۶m�����nl۶m۶��:��9�|���z���~Ƙ���gM۬C%�RS2
=����XX��85]r7��YJ���VL���{�ۨ�S���������#l��D�����I���&�
erGkϞ�NN�n%j�8�������2�}�#���چ�RCSˍW0�B��q�b���M�v��q3"\\�{�AT/�̱��^�0y ����_�8�(8U8�뿔�x���M�U�l�Ck��&8���z�*(�����+qg�N��.��tz�y^y����B�D��K� 2"z�ں��+S=��Dʱ��9���:^�٫X�r�@��������eren\]^�$�IǴ� ��a�~R O�z�<�7b4q�C�,Aǳa��0���"V=怃�D׍@�������P�Ln����6��B�����v
�oxm��c�K�w�=)Q�F�Ň�ݲ_�ǻtH5�!�����a�ɇ��o����pO`lW�E4w���3��*�9k����*�|Ky����H�3c5���\��lc���k"
���e�W����5����zu�/ւ�rI��\n2{+��B�u[�.���OA��8$������2~A�M���� �����J�b��?��C9�ՍSm�i�O��O���<���</N�$�j@�21�~��U���B�t&��	��#����� 2]�pB�M:���*M��N\[ن�2'�1�%�-�%>��g�J0���Ov%���O��Z�H����C�C��W%����\5w�['���J%��
I�E�	Q�,�Sm~Z������\д�V�^�.4�C�t}��9�[��e못�?Z�٪0���m(J
�4Ɯ$�+A�l���{"�,*��d�+�꼺�E��1I�{�}�t������8���ʠ=�	�'w|*���k�^�<��1�ښ��(v�fa�3_���%
q�-�p���2�Y7���¥���9�Q��������J!#R���LX��A2A9Vu�Ƶ���v:��C�z� !NR:�����\�F��cj�!K>PW ����i	�W��p�?=�a:��w����j)j(I�p(�ʘp�b;=���[��]���J(��Y;����;F�xF�oACss��V�۟��HM;�}~�u"%��B�)F���T�X3d��9�X&��.�ٺ߶���<�{��]��66 ��QAA?n�hqp,I���
E)%�ؔf��@{�DS���$Gn�D:y_7J]��.���
�\y�S���)���&�7�Vo�Q�{0p�*0"�P76��p�7��%�6��S�S����2�"�Ol�� �dy =J7���{�]v+ǔ�c���UY�pO���׺��I��$��A�~�_5"�??J��n��@�?YK�6w�N뾞e#/�3h�!���6������|:Am��*	�6��ѓe��������-�Z5'�����(�Q�����
	�c�K/a�Aj�v��ā�I�?F�ג5~$T��w�w��nocQ�sF���)gׇ��a&�RߧB�2Y�ɹ7��sYI������k0E���2>	B폒Q���1���f����&Ii�8��
,�p�����c�Q�7s�A���������u�!{IP^]��}!y�h��z�(�0�I�Ǉw4��.��㌯ߛ���V^� Ŷϓ��fC��n�׾��n�*5����Z�����E���o4]�����%�sdS�k�}<�p�d+���>���,���IS`�aD8�0�{f�$ٚ�61��SF�������=���}	��������ͦ���g�Z��%�/BĈB��������7���b8>N�?�74i-;��7Z��b*oo	[ȭ���܃ʚ��z�"r�����F��ر^KE;'�z���>��~���vX������������=>�fA+��6��M�����G��_�a1�q�[�~�(���E1�غ݆�V4&U�G�C?g�S8�-��.�e4����\��m�׉{q�Cm�Y�3�V#�[�/0�*t���8C�ةb��.�0�0�c�`i��R�4t��C��� ���F�냃EM��JBQ��Ƴ�C���c\�@M�Z�ԏD$NEn��$N�� \!��a]C˄i
[�v����������섐�Yǝ����i�^��dq$�!@B���^�jvծ�����! i/����G�iξ}��5���cU~)lq{dq�5���߇�u[�v�-;F�*� ·ُ=��Ds:S��lUK���!5~>p�F���8Q��m�(p���[ԹFjNR:�@$qN����f.q�l�$�mgL��	%u6̈́��1�1Ujzݤ�j�qh��R�,�~@���DP�Z ��;Zq�[T
W}}F�	F"��9��Y������ìQ�H����2�����v��\q����z�E��s��ߔ<�JE�!G�Sp@fq�*�'O��G8�BYnb"�� �t��V&$�az�4DY��1ɨ��e֕D9��OU�
L}u���m��$��%�q�h�������TJ�Q`�S~�Q���8�� s�ޥ#��^�]�dMP����E"�h�/�\�E�p�0$0'-�o ����$�0d�?���g/k0��	�-
�ڌ�pB�KFe��� �K�&�����7���z�[���?�ɴ�nf��>/Qo_V�K��?2��������6>�%9�W=o�6:&� 0�lK�lΠPn����Om[�;
k�Jc��|�W x�w�_�U��>�Y�	5/��
r��T`�ZB�YF��cwK5>I���>�~F���5�p>D�ؙ�����)>�L��)3��q$d�c�Q����v�uٺylk�D�7�$U�]�x�t)��f�������e�9y��H�6��ӳȳ��Z�Sx����8~k6�f���J��H;r����o���e�@;�ޖQy�3�N�/�퍘�(I#��0-J�G<��l�cm�=쿱Ƶ�ml���T�%:x���SH�L>���D\�z`��<�sP����܆�~�{B�K�M��~��}k<a	艢S_T
e�'�y�<
=�����NE�����h0ѧV�'g�J�����9�7��и��6U����}����#���rٹ�LT��h6\�Z�1>�ں�,���J��F:�I����;�&z�텠cb��ȴg!��_�K�/5S�K�O)
��(�-��D՗��E�;[p&�K�N�X��V"\��
N;98�Xj�l�~�V��̟���9 c�F���E���׬�9�;U���)��\("2��W�
Џ�(���]a��]³X!��nEeפE�!W��=}|�]f>�@���fҭ�6����H����i`c�x���b�2 ����gF!~�H�D��b��/D���r�	2��~"=�-�L$�Z��~�����#\7��^���d7Jmv���Kٍ�4~�5φ�M��^�r���(R�K�V�pŒ�Yl�օ�r��P���&����h�Җ�Ƶ�;YS[�h���r��f�P����+u��V��Ȍ��o�:�I�2<��`N8�2)����KwAD����a��>��\ (ROM���H��?�����n�î܍7��F�"9���GO�@���~��9Qʓ�2��4HI�����0��J퐝P)�,"�Fn��J*I�],W�'l<�c�g�U�j4"Ɣ�
i#w�Ly2�v��Gs��C�����C���q��M�o*��PT~����^#\PBT���L�h�Y�2r�*����y�k����Y(sZO�HL�VL,�P\��9��%5�&���6�Yh��El<O���mq�ąs�<R�I�s��8�(f�R%�i!3q>"�}���r=K������Rp�|8�v��p[��$����ڂ���7͍(�"6^>AC��2�He
�h�~(�G��,#U�Z�(o�P�
��v
:�D-\�� �-HL:V�S&��s�p/!�*���7� �����ͣ���iKc��o.�c������X~T�
�4T#����[t�`��.E��cȴ�E�\`Jq���?�#JgqA��CJ��"j4��^-G��<��(A�z�����+��#}w�s����bb����/7B�>����N��0��@q� "��{3�2X�<As醖�OBV��c�ie5,]���m�C=;�0�r��jk]���
������;4��KDO:ݲ�^I��������-V�,+�v�~��
U�0���'���������W��eȈ|<3���͐O8W���n[4g�����$e>���y[�t��l	M5ZؐN�^�~���m�$M�W���@���q�e? #�=���wC���,E���2�mUi{��2�p;���t�l+1)7��D���`	��I�D=˘~og�����kL?zc�D���NS 8e��jt�[ƌ��UvXL�n��	I	Q����s�)!6�Rq{���C���f�\�Buug�i�&+�LkLy�|���K�W�d��xȬ���,X�}߳�;��������8���0���\P5dtȾ�����W��=��XG\��ܪ�ښ�|D��}wkd%E�'��pI�̮�4�6+fL�J$}
��Ep�D���s(q�{�?!X�> <�K^��e���w�½5*�
�[u �i"�ǰ+�0r���9�~A�7X���K�dM�r˝%�A�Z�a��Y��{R�@���0�:�~��%{9+�^%0�ō���锃�g��n�D{m�x:+��ȅ��g���I�9t\�v,��]͠�t���Z��+W`ֵ9��`�ɑ��P����MÏ��	8+0��B���?�~��~/��#�@[��^T[�� �D6� b���#�"F�6kx�H3%�0����)�.U�E��q[K��k�2�#G���1�Q�x�Z/��5)_��kv��n�����H'8�F�ȼ`�	��<����A/��اƄn�)�2 #��>�ͨ�uX��qЄ�'y�ȡ:Ǧ[��`:��ZNNN^����L��+6<��G�}l!Lb���_!m{��k�_�%�q���D�IL�egd���b����%(`75��ޝ��I��q����w��&䁫��~�&�3�4�Ujme�U��a�;9Ŏ�XR,���BѬ�o"����&:�#���ߊ��]a�&���we�m:��.r2���7�����>��Ek:�3p�J��?c6]�#h<e��~�M�ꡌ� ��Oք��ŗ��8�qG�	�<)�!q�@On25��|5t�\���.4��-��eߕ-n��L����u_ݍ�_���i�(U���(tm�}��,�l��En5%�.B��£���u�6_���X�� RPoJG
�{�jm��Rl��'�0��?���iY��5qh�}��סZ��8E]S��Z�i�����OP{�+�ɀ�#��K�n���"����X7�\�)�����\���pzU��jx�4�����Fr�7d,l7�ۨ�I���KV�i+�J�2fRJ"�����þ���g����!d!O�Gc+�}*N���\ߪNs�2��A�FJYR08�A�>5M+z8;�5�ѫ��\�H����]�1�8��<�j,u�
3q(���@�[7n0�E8@&"�K�Y�(��r��ZL1!�n�=�1��T�7G�vK��-�>�9Ũ�T$�BӍ��eF���k�ʤ	W�);�\*+�:M?墳�{��Zik}	�4�����RK�|�8��Vu�r b��̖'�z�lz8��%3<x�R��Q�E��0>�?�)� �$��}2�T��b� �H6���牲��6��?��6��٣u�T��Z��x�5���S�eR�F���m�K��m*��nV���ʷ���G����St�N6���.�ooR�Ҧ<�Sね�`���6>�.���S}Ŧ�ɖ������>Oؗ�u��U�)��&L����t��r,Gϗ��2ݏM�
9�#��jS��#�qi��1��ݑ�1�7c�|�ۍ��U\0[.ۆ����Ώ�&(��]�:��>�j��J�y�7��ns����)���y�D8Y���S�B����������ܭ�I9�y��ixC�t|ZS��:�����i�b�zpU����92HsIp��a{[��)G�L�x,��D*a�j{�l�o����B.70��]�t��n�rX�[�2Ok���'~����yb���R<#�ϋ������\NO�L������=��_
_��3�_�,�-��=�O"�H(�먚/*�ӮUt���|��*�+5TԾK�쟄<��� �L�㳝W����W�ۯ3��>U��`�@�O'�V�L��	�+u�����Q���e���Wb�ǁ��%A,��{�i�� ��x){��6A#	]X�Xf��l��xtb��O�h2�ֹ����?I|ฯ�\���xx�4g= �Bj�M�pb���!q�T����ߍ��Hhs`�� @����f���ZV�����a��p �S�@Z.L��"s��c��UR��$UGYq���jC�t=���͗�V�����ߏ�������(���WWE�qV�V��i�(��.O�����|�1V���޻��ՅxgX�"��C��b\Q�4���L�1��O|�����6h��(1V�&ʄ��ŵI1��B8t�Nƛ8�C-uY�m�$�x���<�Bt���ܷ���Fg1wF�`|�S[=��hU���~�[�C���X�l����CŪeC"Z��,�-���{H�P��ʂF�)�h)����2����p��H�X�޹��m"��A��m$���@�Tq0�.�ųՏ�u?�Au�n-�Q�:Дq8?�Sm�֨�UK�CfT��C@B)��Bv��P����]�~p�KJ���,��J��/!~C��籑�̜�jj���	��@Cc_��u��с�����^������ W|�����t�P������;pR%���Λ�*OV-�+��a�Ϸ���f�3t��e��rk��힀;����\�0L?2YD���Z]�B;���o�#C�s��oo����́�{{Dw/�=o�ޓOW�/�9�k9�������@f�f�?��#���p[нg���l�P��f��m��AH�T��Qq�oh��Hc���F�`	Xp4��;T_G/#�ϡ�f9���$κ*o�.����4��$�3.�2LW"���U�銠�; �i
� z��67�(jD�AHZ�y�:̸Dh�zs.�|����z�ެ���BY:VM�O�GW�}�,;ǃ�ۋ��o� �lDY�˓4�Ϊn��cy��Ԫj(ysEn5�5��~˸d|�L\)S_(_�{��6���=T������0��=L���4x\��\[rqւ��fW/o�1��8r�W��1���������.�[u=�1�Z�p��^�$�`s0�@é����@N�o��LÒ��� i`��n�R@��<� �u���d�;��:�Xz�|p�Jz���LNJ�*���~�5�=� �n'c��$�/�j� �)�@�"S�T�������OVm�NݺS`�.N:P���;[Y�NN2Ƃ��K�ܸ��y�g��PR1��u���\Zc_6g�(�b���~E6�x�,��sw ؝�
L
�/r)��~���A��i��*���y���4����uCy-q���P=�ƴpr��+jF��)p�%����4�P9<�C+��lrM���r&�'�R�3�C�)K�6ڙ����i��[|m��"�o�#jh0����玦�o�cl��X����$0������y.��G4�td-Z�MK��̙>�6�u:�[�
C�L"т7��I�)vVm��%���}�&#��+r5F���K-��z����+];��H��D�Ę���b�H�t ߽�{{{��y������3U:<A��-�u�ю�����t�E�ʥP����tx�eZ�m�6N1�	� ��Dڒ��v���e�B���y'�y����A���?w�Ҳzf���^҆�p��Ѱ.�tvn.�i3��Ϊ��6]���| ��D��2m�Z�|�E�;�0$Gt�Ŧ����]�$�\�pK�!woX��ߐ9{��WznH����R��^B]ŵ�dq
����\��<	�̃�p�X�J޿NYDR�;�UzR9S�h�G����#�1ɮB���a����ԥe��`�_��Aן�\��}gi��RlTTB��ɲ��p���Hḅ�U�u����yu:8�M�u<2����;}��3��c��0��	>�on�T⹍��R���v���Ѱ����I
�<���)�b��ꥲgK%�搑@����!�*�͵�rE(f�rh��2ϰ ]�P.P�f�e>�/LS\a�6ٴ?7��#_ �(��+�d�;p�*�3@�75�1�t���Zh�vɷJ��P�v�s����� W,�E۬������U�I�f{db#CA��[�]��71ڠ���r��>HJ˖4l���Q:���J����;+�}���+��"�=�<r�s���������X���r\�1|�e/z#z��mDkp��9dT�t��K>ی�ڠ���
2�����{3���������kI������㛳��!��{��c (�ֱ�Xo/�Sf~��>�*��N���B�[`C�U=赑q�՚���t3!jpk�������U#굾��0�B<qw:�ƺ/�p�?��}�g>�]�����}����]w�S�nr��^���Mҋ�b���
$��hz�{^�l��;<t�Xɋ�VB|�GMQ�\j�kV�H�-,��7��`��pj���:�a��y|Dxi�y��y�j?�ǠPx�QH�/^)ƖZ�0uD`/upwog@o
O�+d�)��`(]�z�aU۷x���Q��]0���X�3"�]�P�/��i���:~p#�!����l�����\�w�����ѩ&��[f�"e��j��$��-�����P��T *l��Rl��sSJ�)L3�4�hM���>��L��N���m�i�^nqc\ŜRDxӷI��s�0��mhT�72h�(����^Sy�A��U���l}{�nh����k�&�Y��
by#��VȢ�ak�q|���ZW�f �[�i�μ3�܂�?�⬶��<y�C��́�C�M�v�%3�1|������{�����b=�%.$�b�LpHl�r��x��z{Гg�R֡��L�Z�%�ap�	�tNv!�*�q�ui�S�#3ן��h�Kp�ndE�3U�9O�]ɥQpײ�j�w0�xy �p�G�'�$	۞�c\<���s����E㎻v�cmB㕀�0��I�}6%����+{��@��_)��Wu{����>Sޝ��َ��Rd�9�j��U^�%�PZ�B���@�^�P���e��<v́�v��R�����>Ї#�RO$��W���22�7?�@���������ҼF�H���>]pH�J�l~Ł���(b_����0��]�����2�l�����#�H�����-_�S���72�_,p�w>�ջ��n�o ���i��ʓ����A���2�wݷ��҇�9mU�?�[���s5��"��i��](i����*I��ፔR��~w������w��T��{i�9���4���O{���r�	YXP�,�y��������<퀶���Ԏ����o�A�G�u��w:�0�j��.N��\g�ѽr>�ZVy�W*�v�W|^t��2<m���ݾ��Dl�kh��_Rɔk���
tP��)� \�+[��i����3���b�1*�	M�z���	AҢ�U�@�YWX���;���	H�f��T�O����!C�[|y�
x6�8��4Ұ?����<�KsTl����KQ���Iqᣕ�S�ְL��$��<���ٴ<I�aIH���C�T���~I�+A5�\Vr0���$�HqÂے�0+�!�sUK���LDHw��O��p�m�H���=�����k�+!y&���w���\D����V֌:MM��%`��t���}D�'�O:�`�e�RӬ|��{}����e{hC��=e�lO��<^��I�8-��nx�����{ �*c�1���or��;\�n�(H5B�c�W��>쿻 ��t���G��R4��/�P�;���=��Ӗ�RLe6���ci�2�%��W���0e�2���5aZ$��*�.W����b�ߟWk�/��3�[yݥ{�X�"x�B�=Ӌ�<G��U�Q�Z�گ��>+�����by�(�v"�9NNN�6+��(B�,bnca�}�&ra{-��B����|�Ο�>;�&{��M~�q�BL3L����w>�<qr���\��>=�\1�<u�{��b-�$6���8��tA�I��%F�0癧��Ŝh[e�K����U���S�;V����R��֩�X�Mk�'~�k��.�d��q���Z��5�K��H��ҵg²�g:���R���\P�[{����p#�,'ãyV���W6�o����D�?�E_]�|ٲ�W��v��O��`T���_VM��7������#��Yp����d24�*��_2�Ӧir�d���ѯ'�r��uۭ ��D�ٗB��|��KH���c������K[wQ it�)*��(���	/яDv�'�5�c|�xO�.��9Y�B� ����$��g��%���f����B�
#N�W�V�|oa8���O�[�W�����o�6�1��;r��$3�\T��w2�zq� u�@|�]U�v�ZP��w]3W����c�:�I������(�#�H�ϕd� �I�`��85|
�+@�j���9�;?�4#�������$m+�_�#�tX�y�{i�������*�3Z��B0��l�2��TՓXK�����W��%Y%J�b�E�N���^3�`�I ,w�N�׃��Yݱ(/7yj������5d�,~u��d���Gv���A�o�,�ִ����7j��I���m�&��)�a7�g^�!���g�k˺�a��z�w���Z$G�9c���%'5�,2�5TT�7��>��T��-JCh�b�}�fے��B��̾W`횝eʝaωD� C_FT�me�ҖA��@������ߥ��[lnv,���ۅ:�m^pL<����}OC�&�E:u�i�8�����!dBc	;C�F�!�f`�"	�T9��(�t���_��@k��m�>�ѥ�'_�o�l}����e�3'kTS7�D���;�)@�/3��C��.e��\�9.���+b�3e�#y��2�yA��%�^�r����;T5��FU6D%�p)������<A���B�RaU��)��9�����r㒁��u�>-N��/�OQCr��������)�� �vW�A��ؒy�y��'��)mr6Nk){�P?i���H���\� z	k4d=����\w�x��r��@�8c�K�aw��:Ҏڽ��P"/�������>kY(�F��{���nA�#�ae�q��k��"�}p��w�`�p����R[I�IS~p��2���+���T[��N�bF12Xw�:�2np�eIV⤹��R܇S�Tu�d2J������Nq��|��Iyz�=h��9�B�y����p�XM��d�뱚(� ��X&�����.���-S֫�@w�50�Gg	��kT�䫉f���G�'cPV����l��y&���0J@F�'GU��zGYJB�]�����Nc-���x�ό�}��KK}��}����7����-�b0&ly��4������r"�Ұ~�����⎹h�xa��Mn��<���r�E��TO2��58\�lL��e��
Qó=B>�;�B���g���׫�7����`T�!AJ�"���'���,u��5�_jjLi�n�׆>�z5m_�M�����,��h�dč�S���h��:F����ѴN�K���72Ƅ[�g�^�+��%��.꘷g�����&_�i���[�ߏ�����xb{�Ս��]���a�V잩����Y*r��$���c�[up�&�GY��02uYG,	CF�U����d��=��J���a���=CWc��ߐ��&E/�?�I,w^\5��ޱ�a�Lıx<��M��Ie��S�F>��ݹ&8S��f�C�7�LPO1%�O��>/w5�	������J�#c���q���nF���@��5� �o�|	���שK��N&��h%0�E�y �<+�x�*4@��(w	�<�>ku��������dlTa5?��H.x"�(��x���߷���Lv7�2d��ePCm�\�#����ɠ�Zj=2�x�V�0F��	sp��Qt茁JrMR�jKY��*cbm���T��_�X:F��X8COO��"
Υ��K1�d�q�N��ʆ_�ʕ˛�]��4��+XI�1�ꈊa�K�
p4�G׸o޽D���q�����xug7y�{X���̀�dHUǗ[m����'O/�-���+��)����5 �ɸqi�x|h���O���2��l��;�!ɥ�R,��4�������׺禀���gS�w��^ V3A��K�v:PX�i���π�(��y�@'���g�QXwh`���r���s5d�aZ��#�}&��˴������U�ċ��yq	�:�r�l��u{����{a!Zn�1B�ae�I��;�~����ӧ|�6ݕ���fk�2�;��.�eb-bC���˾��������m���ϧ5�ݿ�Lj������ J�9�3#���Q�MI���M�O��e��7*=_��� |^�QF��E�B��������mt�T��Sb� ��h�y+���:AN��Q�z�&�l)�T���[�^J�A�ҡ�1��,*����ŷ�Z�z\��5���Y��A&Xyn2t!�4���
���!���_��*,� ���d8��y�&���t3�"�hġK8z(���m+�p�-�bp�Ƞ��-�x�^b�k��AnC���X�+)��$\)�q`��Yb�4I�w��2$�`�`���vɥ�^apL�$�2�T�4�/�82�I����uL��l�HB.ս/���gZ?�E�r������HЙ[k�����Hˡ-�)T\h-�ɒ���q�[��&�ހ&Hw�ZQ���̌��4��4��&���m���%w�t�i�!J���"�\v�q�J�r�T�Z~��	?���~xi$�%~mfb�w\%V�))Q+�+Sq�����;�F�}6��䅅lo����ݗ��>˚r[�.g1��޿���H��B2�Sl�sq��7U%��R�h�J�=O?娨����ϐlP૑���-e�����S����)���~��/��%��_�z\%yqp�J:�Z(N�[�'J<���G���1��J<���'�K������d
FJ`�U?�RQVc�^��W�@q�{�8W�/��P�A�au�ڃ<��#ߐ���ecb�V���v`�6r����A'Š��sk�S>L|�'�T���8�'&��H��4O���ӓ+�~*��ˣ���������ޞ�2������ ���qY��&���(�E1��iS6�+��,����?}@kza݀,�{˵D7�֞y����2���ջ�$%D�!���N���5޼�ZnL�l�r�`=�͟��&E?���;�e�İ�/r����b�d���R�CY$�GNS7
V���R\��U��a��^N�F������&"���@q� �>L@��0Td��E����q��@v�F�Y�T0�����&�ʶ��6��,�fxgI�I#�g�����4-�d�%?~^�1
I�5���	^�贇;:���rL<Ԥ#����g�����Iyɰ��eڀk�u�.,~,������H��/��re��QN��:�S�$V.ɰq�]�d���D;�\��m�V㎚�I;*v4 D�[� ��"�4� y!+�0U0p��޸��f9�Qf�)kr�)�h�J˸�t l`U�]�%:"Fp'J�u mBy�^,i��B��k��J"�t\���Y`R�Y�)ص�c�/��`֚��"Y'�&Ө�!c	yq6~�@q����(ጵ�a�H'x��z�{��[�#`(�Z��L��
׻���0#��uB(�\��J�W�E%�����T�6�3Do������΢��rdi���nB��]��aU��>�������Q������J���_�M�t�<KR�6��gnZ.q{��X��>~m{�ɽvS�z4��8��b8)d�?�����xy�۔�KH)B��EZ<#~���Rt��2��N~w	�ں��:xP���m����^P���s�����a��>Or��H�r�'�Ŵs)�����լ@
ݺ8��gOG�n!����33�|6�=�f����R~d�`E=��W�)0O�qI�A%?]n�h��+1Y��ς�{��� �T(���1ІT�L�e�e�r��(bd�K��b���ANK�J���^���q�N��Y9z�#�����)�b�e=�]�P�X�19S��0瓇��6|��ų�m��%K�&'7��V�ڏ� 	�?�f���޻�+'�=�J��}�'6��#�	��Q��ju�9O�h�۫�ɬ[���*w����-
���/����'L���Ģ��Iw���/��*��SR�9f(�.é���JM,�)���!�p�,ixS9X���x��>�m���Fb��z���H��F�.��~��Ļ����)}�����m->�E�t�"�*ep
-�Ku�9�vmQT�+u � ̽w��W�������8��~����o���ަu��<WX�a4��>A��7�I�]Ϫ&���^X���oOHW�T�4�`��G�jjIG�d�ôI�8ݾS�[��twJ��On�h I�bQh?{ܼr�>5�����z���|��q�2�?��������#G��|Y6�n���j6��.��!e�7�'�J
�0L�#�3)S^�;Ù����޽����{ŦiN��9FzP!2j��^�[����b��_;��d�3���7��K2Z,���v�0�=��Z��6���7�$��=���/	Q�wP|lԶk�&^!�<LD2	��>�%�|Ey��Ѱ��{<����`R�֖��r<��Av�G������Fz�	�+�{��ǜ�F��CW¹��U6�j�����+��H�I�G��1�%������[�>����l�KFJGB�	;Ѳ����ʖ<7�4�iDյ�AިT/Q�8�V��t��ԯJkN����Y�rX悁�$�4����O���&�ٜ��[��>�}H	�N�Kb�Q|��>ꄝ�d�$���2��Wy�'�N� V'UC#LB��K�N�|�Fv9��"��{���i�q�,b�\CO�E,���<�YM�(�|�g�#�o�)ڃǄ&�:DXx��?-!��P
�@F[��ٻ@���h���!�#n6��Z��e�I���j̐�JͰG^�qv޾]W����*7��b!� ��,�"ڿ�o��r���]�|��C��LX����qb7I�K�������|rae�0; n��b��Z�W�0j*����ϻ�nQr��"V虁-��>) G���9���T�z����]�>{/��A�@j�����iRT3��t%�d~��~](�Z�ct�L�������j�|#L�|�����\�x��4�E��|op�7����qMe�5S�l���I�����1פE�t�����T��w��D�r���¿)0M�����cK�\k.�umU�EG�j�]�c`�K�O7��b��ٶ�d�k�]3aΧ.��7Jvy����=��m;�Д���E��*�V���Z��t�I��Y=|�7��u�N��1T��d�,I�RE�Te���c��0cv�Z�&v��V�fr�S�ua"����i;	�.R�Y���A&�0G�Y���jT>�?*܇�Db����( �<XGT�����|{��$:�g�09_� � �A2V/�A���(�tq��� f��E6��ۑ�?��u�0��H��H	~
w���>Q�;�g��匕{�X��mT^$\�[~l�yo�[�`���	��'��U�f�؊k��M����>�Wd�R��G�)+�~D�V�оBZc�R��TZV�*��#�'����R�[*���yN/�VR�#���4��Q�*���qO��S!�ǋi% Y����,���G�'��.�z�y��E��%�Xv�|I��5�����T��G�=.�I��6�Y<��R1��5�'�U�_� ���	�:W
��D����°ˬ�7(��Ʃ;��)�?<}s&���ƶm<��llll۶�ll۶m۶m|{��0U�g�9�=ݕ��@���A/�2�dO�غ�9I���
�[���c{5�)���):�.��reW_��eTkY�>��T�e�R M����8�S��� F�I��L�Ꟶ����?ׂ� �{g�&dQfE��e`�K	 S��%��=���\�:ѷίh,̳�9oλUg7�`<�8�*��>���ɻ�P�� 0f5�'�~x����++�![v�<0`��u�'����	�u���us��W[S��i���<��#�8*�!�9{4>b�v����P�k��1��Ո��]�Q�}�v��q�E-xF)�L>.3�չ0Oَ��k�2o�҄��9CN�ޛYߌTń�Z������[i��*$]����s���_fu6k�%j ���uɩ>�fm8�kh�[�ߎS��<�:��˞s��SD�I���%>�.��T����u��˩9��Q�$`�ʉK�"�uP^Z¡�7��7A�����=já�M�Dq�f��mJ~���ON��D��D]�\�-(OxD{���54�L���'n�qn�]�r��|�:��A���3_�6{��d"H���SW=2E	�ߙ��v[�Q��ө��AQ6�$7�Z5״-�D�nx6��:�������>��Ƚ�u�Liy��g�*"�et~��F��;A���5����<<g�֥��� }� :A�4g��/%����w����3�Д��Q.5G��c	�>va`�C�#o�2��)%��=��e��}6��L��د�E�x,_���-�Un��#GY�j��i�*��ڽi'u�4�E踪<��T����ܣ^�o�\��/���98���Y3]Np�ز�V�,����f�Wߎ�AoR�T� n��-��C�Ұ�O�K�R�zg-�0N�-^Q緯���+0�Z��Y��F���3����j+<ѫ��WE�zL1$b!�GϽΨk:���yR%tA���?x�?k�
��^\^}ѹ@��W�*��,d3Ƀ��Z����P:�Ab`i�3%%��m���������DVN���sol���ddw��νN���&:r"�f����1�oԥ�^�*&�}Y���9O��@C� !/(ݰaJ��"d�g����oF�K�Ԃ�����*�[�(���%���D�����BSuW��5�\_��EF#��J�ܒ扯%�b!���o�Ӌ2�>2CRa��C�� ^���^�`�\��b4�Aǵ�^^N߅h8���-���u������]n���eics��:ih�T5�߂ɔ7*3�:Lxb�^�X���C�=�D��-x�a�(N�$N��`S��[��D�e��|��`G[��q�Z9ϔC�� �ʟj`��J��(DE��r�Y}9js��	!��xr�F�xuh�oP?��8+�[�Ǌj��@��w[1�Xsb�@�:�`4�B9�QU}��g���&�´������q��fo��{�iR���f�*Y/���.�4����)F'�}��Qb�{P^�f��eW��R�����Z�v��T��%��D��,ͪ\��Ul��
[G��	�]S�Gb�:�_M��	�OB�mXN�g��5�^��h"����0�5�/�B�K^�5aA,��U���� @2k��=��>�:�&f�o����p�+�/ UXŞ��e���&��/Ҥ�p�$K�[�b	���E>RC��ް^�Dy�z
P��YHn��uQ�?j3I�"
�i�+�	�~�_�yBY��,�|���~��D?����5g�˩�t��f��l�"�`��$��<�<�
��5��x���!���F�1㺗����C��-=C-=_��߶?#���ߗ�٩�p@��w�lY
장˥Qk!ܮ�Sǟ�9��A��:i#ߏg/]'��߆���צ]
����8����s�ۏ� �	����)�E��4Qm�P�
ӗ�ʼ[������}���'�:�����e\�C�gs`�_K-�
7y<��O��\����Yw [��Q[9�{��P��Zx�d�;#7p?{���wa�K��C��zߑ��e�i�����oE�?c��B�.PUy����۔ ׆�T�T����p_]�PA�ab�^�s�a�J����v�L�0���.�̓�>�p"�ս�%��	�d4V/*<v��R#��$F0�ό�ӄ]x:�f�XS�����M�sJ|N��U-!�����}
2��t�T��F��5�Y qS�#ްL6r-��Ԓ��idD��z��"U���m�ѷv&�ӣ\�a����u�����)j�����mzDn&wsƷ��F����b�=>�RQ�BƇ�%4�[�=���Em$,�m�>;+l�@����9���O�t��k�Pm�O=�J>�"�"�>e��8�����7P��&������JFv(����Qđ���T!Y��خ3��T�������Œ�����Tc;z��v�s��c��礰��Ϛ��X��然CUWy���:Vt��V�BB�}�p�8)$��սT�(�w�a�(܆�߫�4�$Vc�h�"ṿ�	Ã�y߀{T]��SW8�Lp��df����#�@���+;�Y����x�����vJ/G�x�p��>4	�

���ƯS����Z����w�o���aY Ty�x�x�d%�;+%�;��<�b�i����tя���?���F���z��������
I��87��Z�M��w,=�د�Lɶq~A��RH��y9�Cu`�Ex�!��,�?��D��T��2-K�z墘��EN��)t��q��r<���پx��_�fu��s�� �J��fL���P�ڎ���u�"O�����o��j���t	%|�ar��u������}�� �Fm蘳������=o��!\T�RaeU���՘.æ�U3�L�s���r�![B^�����s�p[�?�8I��\���gԪє
ѩ��n:�^k�ņ�{O��b�nz��Q/�'�s��_H9-_��0�0���]��ՠ4�S�t�zp� ρ�z�\0�=��"�����P���������2����&~�^C#�a�M��
��u+��JV/��RfFP�����Ӗ�@��RC�zX u�:�.ՠz}���#�(�,N6�{�����O�w۫���hHY�{J&�/�6��7L��Z�Z�8�)�Ŏ�nil�� юD��5�u+�\��T�NA����7������Ţm���q��a�{�H��m��.ͣ8ޒGa�7?��ә�|
Ek�Dt����D3JQ���]�r��m�M-��</L�|�f�T�~�d��n��ZW�����5���h�ovQ�0u��e�b�`�H ���IԳ/��[����'�����h�*�ir<�u	%�����3���"3j���	87�f���h�к��Q�EI}>R'�l��K��$LN*��	j�P�L�j�d�4��_���ld�3W��1�|�	��ez����͟��Ds�Qn,�墔����$�rIn�#�+��բ�)�"��X�=��L���l�aT�R��Ƙ�a�֨@�����ևnD�cϿ?��,��I㩓�A�*Us[F>�9�6�ܞ�3���������G�� I��Y���~
��YŜY.)&E�DdfU���Օ���7v?�����{<�		'ũ��ݓ�0;�������9��e�}l.�3��O�	1g�v����'L�Uhnr��yCr4�R&S6Ne�xPB��34k��'Ǧ�K��U��Қ��^�fF�2o�ʠ�H����A=	IV�g� �C_���F�F�oה��ݫ�����g�����e=���	4 eD�`a=�r�"h�O[�]�L^$ ����pmvlZ���,>;�.��w����6t�Ywb���&�<^�:P��23�o	�3�>�D\�]��E6�,QR'K�)V��i�ϐ���_��A�^��c���ӄ�������
j��ր�F|�`P�G)E�J�k���$p2wߧ����+�b�����#�}��l��
}�~���0��ߋ���	P���F|�Xn��#}(��2���$��@����ѨV��怇
�e�\O3��E�V�a��xh����nPU x�9��)���gcˇB;m`��QӿA�J;!,2�O5N��2�y�g��#NfD+;C"_��S����nc��#�鹲������Z��Vf�n��N-%�H��=\�T?�U�V��{*��������5���K�ű{z?}�6`�ܬ8�%eY-3�|��Ò�x>W����[�M�Z�!�bu�&�7��谆��;�P����$c�����iI�@���û�������h���*ӈ�*t��z%c�O�>��I�-��Ϯ:�)	�<�����M��$
�֦�;g�����G���[J��5����.7�Jd���ť=3�{�OMh���t���D��D{ㆶFU�E[T<p	����
��^?�u��s�wʬ����O�)����`nW;G���<�*)F5M ��i+�<��8c
������G�9F��L��㾏Бa�|bf�#�3��(U��	c�mig�L%E+��U�w|($������Ƒ�$� d'�9��֑OM2���
��+�]���zܵ��}H��I�:7��Mٳ�c�D���$�[1�{���x��a5��+��ȫ�(�R�D"�6�M��ln]k|�:�۽�l���CQ��E�K����ם\.�����i���2Q�=&�D!F��v�':���*E�<��o��@Ԟ@M�$K,҆k��k�h֘�ڏc��ID���8����&0w�P8LqV6уg5�[!�N.�N�%`&����y��Dσ;��ƈe�X3,y��@(94��
5V���4X��4H�����bJN]��s�+��4��c�+���8�1�Zz>s
<~��Ce������Q�a�`�������;ɩ!���hx�΁�H�mg�xk�P�d=b.SL��-"�~؆�ϙ̳w�ȗ�g��O8;݂��ȹ���7=&hߡ�$�����S���Ps�?.��[���I�#<�a����p��q����eGHi���?�����4�em��	W��!�)�^]�)#������ԓ��ʆ�)�_Z֬m�=���Xm����箖�)�멁�����#*S}	�	��Wu�M���gx}�s��� �I~�r�'���S/�n@���@��a���/W��� �����@�Oӛ���2ۻh�OG�JD�������x:�{�+�P�%���9�*uMmCg�'�ӽ$�њ�N��#�������-Q3Xl���?�Q�s�_�A�9�W���w�v�4�Fi$N��S\�g3A$�,�-����¥�*�	;�E��厬����U�1�3�uk>�Y��yZU�'���%��3|Rk�S�;F6ψ�Z�K��SZ�b֫�8c3=��-����
j������`���&���{|?P�ZnI�_�$����TZ`����gh���V(�;ւ��8��Of�Q����VmZU�G&a�ZC�<�|�2�i4P`��yM�~�C�^mJaw-��t��aB~1���+r?z��jy� � �j7Q^t;�^��pkE@R�[���}aHm��J�XIJj���0�I'�VV��QE:�+��́��Y[��{�]��i�����B���Ɩ�0�A瓸��T���+�R5��@v5�T����5�!#�S�#�Y�H�eQ�Ο��z\�b�S&���ڳ�[�}0\�^G��p"a��m�dB��$��$J��b���� �m��\}*rZ9yL�S6�p��rc��V�T_��;y���֨!���P<k7 � ˙FT�t=PF�Xj����EY�J�t���-m��� -g~��;h���C�-����'t:\�
b�j���+�{/� !����a�;u�[_�-�}3Q��6W���w4pV8[�'Qs>7t��\Ϝ[�Eێ5m?���,�Xd��3�o��lo��%ۙ�,+��m*����s�����z|_�o궐)y�³|�
E���"��1*�	r��E��bsa+K���r�����C?����jY!�N��B?[F��.%�X�Y��6nW�[�K�Ⱥ�..�h}z��}ߤp{7U߱BI!?��d�O�t ZX���!�㺼fI��{N&�P���~���������k���d����iw2snǣJbҠ�ֱ^�x�L��e����;"�J[Y�ػc�-Rʈ��,l��@g��(�Ri���`���{���o��-�*
7�"��j��W����T��+?=�UCݺ%�� @D������Ꝝ���׷�L�-��r��u�f�G߫$�Q���%!&.�� ��z���F���ˏx���A���E���	�V��G���0���)-75k���v�l��9���F>�[A�f�o).F�\& �[6�!�X����v�;�5*�� �z��}�aSo�߭ {�r`�j4aE�(,� `?�o~���[�&�p�:�H�L�O�$�䇊�a����x��25�ilw�N:P|�����~!䪅U�^�6�e��ON�:��8{ ��ʤ��CP�NA�R8Us�"�E%/�Q�,ٔJO,��Q��>�����2n]}�`��<�2@Hj���&X��~~NΓe�6�Im�������ye%E}Úp ���"�1y�x ���3�yM$
X$�)�[go�wV��>)�JN&����Dd��_��o�~Sp�(���z_m�����mw�	�QP��}�o�Q-6����뢗��EZ)A!;	���xn��ZR7i�قe��+N���gQ��i���XӤO������ۇ'q� �5C�28�T6"i���!(G����E�%ѫ�h2[3HZ6GΥ0���K"����I�&xD�.���1��Z7���	��=ov�uFʺ�j;���.m���G�^�-�hșA����Y:����Q�X)��q/���I���]��{�����6�rD�X���A��%�Cd;�p�Օ�0��9I8ԛ�+WN\Y���C+��s���%�˱�>@U��)��Y�n'��l��-�KVq��Q�^�UD#���B�	��%�^<��ϻ��)n�f�^%H�:�l���aٯ�?G�Ŗ��e��6���TW]��J]Q19)���>���+P�sd��ʔB�{���~C�iR�`"f��_X>���-�.�o��<�4�����v|����v�l���BD^�� :{Vj�����3>{�w�������s��s��*p�x���%䗤�럧7,3�{e7��0<�5H�~�©��T��9�1��\�y�����8�V�{��0��G�W `]���D�a�'��<~ݓ�$��2n�4�ah� <�m'{�F^t�s��L����s�]l����<d���~>��apt��Ѧ����n�tr��n3�k,)�f4yh��&$�Y�@l	`<�JM��g�O�����G.�\��P�����jrrk]s
4Fav��Q��2����>�ۍ��������ٵ|Ur,����uc�2�ZƂE������N�ƙR����p�F5]���94W�~c�9�hW���/B.N�7��N�}4��~�Z�`Ӏ^M�Zv����Ow7Lɼ�q�R�&Ҳ!��&�:P2�R3�u��dTw�P�hT� [h�i4� ���*l�M���3{~	�آ"p^���i�?f%1*�2�>Y���M�t�å�Y���|3�g�Uˢ�y��(?���qy2!�b;n:QPd�l	��Jl�V�^�',9�0�0��FaIhT@1;	��o�S������Ch�ӏ�r>8��G��CƂAH��m�>�f�n��(�Oa�~!�'��
���ʿbM��!�Ny���e��q�f�����W�*��>�cϳ����p�ڇ%�[4�S�fy"��wU�_Dg����t������X���G��q�;���_3�lp{C��7=ɨ�43���é�{-6�0͊�eN�o�`�0Wg��:�q-������|P��i{�"aT^	.QHV9�Xjv�~�����H)Ԇ����ӻ������ok� ��|�4���ȚΈ�t�Y���!'hY|�����_�yɂ B;�hA�P��ά�B��?ꥪuT�9841oi4̩4@��3�/`��Ǉu��&�ϛl�njۚ�ӳ��Dw��^�T�z�HN#ܩ�#X��D�r��
׮��c��$}U~�V�5g=
��Ѡ�7}|k��Hi�
}�<�����[ĵj 	V��	gr��3��k�5���-<�?�d*C'���������*����=5o������]L�R���:ȳ@x�����<���K�b�gn�qj�_����_=�N��_K~N�6{|3&��h ���?��+����k���8���噷|$L|:(�L�I�b�V�G8���B˓�̼�K�c��#)(����ed#�}�k��P�s������
������h��gG~aA��>؎��J��\H�)w�Z��E�/{��-�@��T0�"0�X5���pK�B�;���m/ݨ�S�T|]�$��`�Zh���!�J��+S��l��XS�d2y�M������E�t)��zs�K�J.��¸߅e�rqX��	�����#9|�@�v[HW�N��>J�1mV-�PD�O��O6D��,H�,v��?�Hi2���)�(��\�V��r�.E��0CL� �ɾpdl`�|�5�yˣ��(��3I�&o�z^�"���JF[�T��V�6�9�U��셻�HH"q��û��YM�{���?��fo^�U�-�T.�I%B�-(Ǟm-'V8}�x`��f�bs�)�:�-�
�
����i��Pkb��t0MY�������+jԁwj����^������&ީ$K�Q��q��hp�����燨4}��읏�v�#oV�9+o�3�Mo�/������״�	(�wӚ��{��	Z�.Y�t�{�L�.L��Yh����y�Q���d²�3��ENDA��F��T��ȇ!����ĳe��L��yV�h�eT� ���k����P���k�C���I����g4�n"�	?T�.��q�p&!��h��O��ُ+�_�Y4B��Q����ĺ~����NF�K�P�0�$�TR/~u�F��W�r��)�K���"��C~�y�!*c�őցG��z��]����G��O�d�`��j�H�����(��Z��=�ZE��D��Uc�AL���IϨ���Apʶ�{��������P�Sdq��K\d�ԴP���,⫁L����絘�H[ߚ����-EKmw� ?#��ȵM�2k�0-u�i�^3Bf�JY~��3�P������<Y�V[�}��u��XP� NM�P�ku�->	{z�Y�2$3�v�r�P9��r)�f dq���]yĂ��|?��F � G���J�7O"8�_H#(e,',��yF��/a�m�m��YH�܀_x!A����\��uuG���os�ѬQW$�s�H"��mW��6܎�SU�j���ޏ�X�T�%���RL�B�mjtߞÀ�m�QJ��5�2'�<6��e26v��?%�+�
L��D���3����?ļ�pyiu�~Q�D���@p��`u�}����;A�<2Lq�� �>_�TZ^O��9��Y�xTQ�dK"B��I1y���J%äa̲�;D���O�8�
'6�F"5�z�L�;O�.��)A�pt ��	��ٙu���f�uuQ*P�����#���1�l����+�J��6�<�qr287$R��v�2p2{?_/D���!�9+���{V�v}�C���4�ܢ���^�� =�Y��U���t��zM��kd�>�E��1m:���a0Is��2ݦ��Qq��%@���\�!���"Ϋ29�G8�b�mbc�..���~�y����}��6C�M���>uڂ-����a��k�S��,�����muu���0�I{� &�d�u\�2�ZY��nQe�+�LE������ɡ�2E��F�T��b�c�%`����KМjKb�����������YZ�1D�C�z�Z8�V�����'�C�����o��_�S}��6���]�p��d:�Lv1O���"���|ABĠ���Ĺ�0�'�'C�z���f�)x��D.E���=s_:���k�M�5�8.�W��H�P�E�������~N������7A�{~��i�!�1����#�a����󷮐 ���-�|S)=���2�w�3�w�ܝ���*�LhE�f�q�H�.�Gj���+���TKLq�Z�^`�]�S���҄ N���yf잻���*�QPa)�h$M�9�ձGXɨ>�_�(?���Ca������e`ԣ_�$!�
u�]~_R^�����������G�Z�$�O��`�DǛ4Ht,���ل,l��Ɩ��\<=��f߹
$��x
KE+@�R��j %��ъ'D���m]�u,�LP&�'N��F��.S��Q�Zxħ�I��Oֻ�!%\�9a��1��
IF-����,�u��P��jɖ,�\��X�7��0ssKuuC	hA˓��0�Q��%����)a!N�_�騢;/�=i��\��R!rIc.��(�B�n��,--�n<wp�>/7U�ؚ�z�ؙ?p�}r���[z�ۚe��v~��$d�.�R�u��I���QTJմ�j7��Nk׏���g+������k���
�A�Z���Z|9h̹��4;:��L�Ϟ�..6(�
21RӺ�t?�r�5O6�Lm<}ɞ̑�����A������>����,M�t�����R!X[qz�V�GZ�B{�WOg*'fn��|��U�7p�RB���Mt
A�
�*�؝v�p`P�w�LJ>S�!�rW�?����������M���L�Ā�|M~{28��?��βo�yeG>�����"D��W��X����_pj�ᅳ&i��R����V!��S$ (�ʮQ�	�--(n{i��#Y����{����/�I'�H1��1#�ukj��H���)�Bj���Gz�O�TB(�� ��f�KH���m�<��}'�	������?\�'d�V>�a��O��.	�d_��"j�9k{��;!i����W��5Q��J��q�����8?���u��\�\�$�T&7�8����L�6�G|����]��F�A�*���eQ$��H��C-�����kɾ<�(��+�<+�R)�(��,&)�~�����L^��yߔ-�&��L�oP	Mn�>�_\�)P���Lf��#�SwB<C_z����{�+HI$BU�"�&��_�[�z��!<3��� jnQMY���س�%�g����_L��RH�r%�
�[�7*����R�
��+CK6���5���x��
b�L�y����rZV)$ф'd
�U�����NC��&������WW�AI�S-H^�FI�Ɩ*b���)�R	3��J�=|�A�6��6)M)�c��h�BneHN�B;?Q��$��:5���t\2Rw��bi�\�����)���c��n�#�����9�������VV�>޷_��3yKI�+殱�u�v~�d�W�N�i-�nY:#F������M\	̡E`��w�8���ev7��#�{�@��F0A���4#sztt%JIU(���`��[U��˦e���A��P�E���|���z��|����bÑ[8��vi���w�>��ip����Oq��7��ҋ?"����}b��T�o�2̈��~�-��h��_� �p���娲�I8�VwJ��e-f z��5��A��>�`@�����}����7N����C�2���~��̿����������S
��E�'��p��w��@כp��O�ZL�@�(1Gw6�����"�y����W������2��b�,��X��`v�'Ը ��(���0U����7�����L���Jr�Y�ƿ���0D����b�硘�uOF��)�9��2}��W*q�[Jq�/�XSW'��%ߜ]A��{�N����UL��X,qh�|¡n����%|�vM�{�Ys���{;M+<��0J��X�h���Y�#[�6���&c�����y?��2��Q�`wG�O@]���	�$���&���}JZv6i�V �
��jά�QF�T(��\K]_d�0� ��%Ц���܃�[�u��Wy�?���Eǧ��U��(6�#�u��%�R� *0ւ�`���@Z��<����3EW�n��w�|	zYc���D6ˠh�^�Eؾ�'���#�� 7g���ԏ�.��~N���}�V����u�tp4�!ͦfdz>��:&����o��U��}�K3�����t7�9�B��蝶g*F���aLe��U��~�~�H�E���%K��9AC���C�R�z�<��¤l褊p�$�A����;]/%*0	�,b��q��*��8�N
���e�$�QȴM��w��P$�V�Rɳ�Џr?��ΩK{��uc��I��)��)�C�e�耫�qh��e�6�;k}�F�w���pi��&*��M����=��ģ�߬ԛ?��2h��iÜ����l.F���Z��D�8���+dX��z��1�N������_��ź/zm��WzG]}���_\�_;_�b�=__;W���%	��aiC�g��x���{�r].�ۢ���q�v���<<�3�wGy���a�~�p��+S���|��� �,7�^�����:�h���~EM8NҒr���-�i<v�3&G�V�LF������ޮ�������Xbm�+xH���<P[�7>2�w�=	���߮^ko<dǂ��P�5Z}�7��k�s ��M�/�n�("/�1�$�F����-����O�#�41�7��ݒ-�7�%�|�^NrḠ�+���tbz�#R��s՞��K�@��;��Ojz{C���;C�d�u޿fTh�W����@��x��Y��5Rj�/���$'w�{�j쟻=߾_zf�j:'�.�	��/�ӧ؂��1�Vi��
ih&Ϛ.h�����쓃�9�q��+� I<��*��8���m_������(�%X�����L�ߧ	��!�����}�J��V�	C��sh�MOfθ�3�U���~�ȾW���좭ͼ���I�ρ���8Q�pE8�D%��6��.���g�a��%d�&�%�����Aw���@��p��]���n�����V�,<��-��\r>�Q$��˿3����W/���K�21�r��d�Ytm��� <�i̦��t�(�4����yG~����F���m��S�6I���%��on��p�|�޽��C�߃��tM�,�y���X�Ή!=/?�|�qk�wǗ�7�@�F���ケ�Mǥ�i[�8~5����	�#w�=����r�
@]t���ŉ �ǜA=P�6�?!K�@Zɶ���V,��k�9d�<�~��5���ᮾ�76-pp2s>e����״>�$ȶL��)H&<{XU�(�%����o�*e���dg��L��/�J�$�E��x%5Y����\�ʊ.�곳)�w�����@�|-�	���l������ޖL��R�1d5u��:���<o��c���o�Eסe������x�����!�#�*��Օ��-CZF�������y�#}�+�?\�YʬK�}�z�Є�&/�W���&���L���z
����ơ]���,��%=9k�;�f��[���;���Pz!��:4�~����kM�:Gl��	����)q�N���A�.4@��������Xxͱ��D�ڮ��I� �.�#v�tV7Zq0*��=@}�AƱ�	K5�0�ޟ�5��H��U�M��}���>"��������I�w�)�-���Ѭ�:}�(T�����O�{���CS"����s�vw�����[>� Cq�"''%�m#��,в��\�`���lzC>��������}��O2���|����樨����'�ڂ,���1Aҷ��ə�X���|���C��0��q�?
�rz�GO�i��C灶�a5��8��T��"�Iˏ�8B�%���l�t�9ɳ�I����O���֣������C��>����1������"540��L~p\4,��!�zh6���գJx�"3���Br�?�H�'�EMs�"�gsX]R�h0�A��s�孔�S]�1� yn�����\�*P�2�Xȣ$�����: )]���W�F�ke��������ڐ�a�n=p4��8�$���{�{��8��f� <�Te2<i��(�望m�����cb䖊^����4q��~�}ߠ�T^��,H$�V4=s�����`EF��BB�F.Y��sg�S.�~���2c�x�i����ۍ�	7��a����_��)��W����*���.�k�������<I�IEE�4;�1�V��Jr�Ha���X[&�GK����Y���i#9��.�"��TGa�q��2�y��4p�����K9�0^�b�W�k�V	��@��Rx'FQ���J �K/�*�@J�[W�"��(Y[�9h�hy]�>�{���Y���\¡�����7��i?N�l�!������'�>W���e�a�߰�cf���+�f(�?*�8,�n�C��9y2��5Ղ�%#��U���]p&f��OM^��$������.��;^A����(���9y^���"�F%�ew�0-�$QFcI|����i���R��1�:D��n����(��E�Bx}�ƈ�p��i4�!�c76�s�hҍ�{�l��Ĩ+m����1�s��l�rh@�J@��%bX�3pF��(a$��Y��ݏ����k��O>Ms�C\j����=Z�6Si����&��/��=�!l�u�}}��=u�X?W�
�!eA��5�g[��n��-<>v���G#���VaWI��腸��J���_��?�?�&S�
�b�>�\)l����\Bcnl���y����/���'����/��?_�3j\�� #�A����m��Z8�)��C� ʙ%P�HD�u���Q_��Uqo~�í���&~Db|�E�p5QD1i\b�n�Q��u�/�a��~% ���:����_=�s~ᗫ��K�Qy�w�Z��	1���y���HQk
C�8�.m����ieۅ�ðF���#��\݀�?�ͨ9a�Jh���>6l:~ lx�������x)i}%A�	}���	��
�&`躧F��tb��BW~�˾L�p�r�i�"�
�9W]��w{�p���bR�շ�EC����Z��g�I���p��(U��`#���*[�p� ����?�Lǝ�*��"�GjB�cK��\JJMqZ�:��R�jc�!�'��������k~�kZ�3z����e�g����ޞ��rdqΏ��ԓ��֔k6^R�'�i�*�f�]\]9]�e�Hc�m*����Ξ�l\ۺ���&�y>&'�ع�A�f���"���(���1O�۸���7�@�)T/�=�^&����D��<Ө��@�nOLN�I��8<�e%��|�|������o�Er_s�hlp#�S�ܗ�!�$'ky�H4���
���{�v�|`�t?�:{���1���!l"����f��D'�h�X��)d��k����āb�/��R�Ʒ*Sh���/�[#j��>�(���ԕ��/��/q9���Y5۟"���GCH�+�$�z�=~`)
��z�����7�~ou�Ն� B?�/�{��pT��y�m%����8�"1ɬ�D��	D&w4+�m�A������,/St#��5��6�Ǎ;ѣ)��� G��W��R}�.y;n�=����ڢ59>�U�kD��4��d���'.���=������r�v?y|o!~�[v|"�W�峲O�@��!��tjB���Q������1�5߷�d(!��5���&y]��~r~2���WTT_�{~�9^�9EC����ZZ�H���7c�9�"�4H)^��9'ɚ諫�nGK�k��sb�ֆ�r>�(��3]��u�
����č��T�xL�́�@��Mq�R����{O�z�܊��ȑ�J/���������<�_��hd
���,���s�2�����?�c��T� '��HgLT�,�A������Іh�u�:>O���	�J��p�ψ�X�o6Ts$G{-�]�f�xT�������3�/P�Ӳ�� �=�1>�tבl��Ӈ ���%3���"!2V�JQh�,���?���|$�(yb���ǴYE�l�:���]www	�.wи�K�w� �������s�}؏5�U��5�����@N~���b�ÚA
��T��W���:��*mn�M��Z�mU��_4��֋���� ���O��R��\�
��A�F�3�fa5d���J�fB6̦w,�R�|nh/!|Y��~�*��M�n`�����Xn݁Ou�J�p����)�n�{���#�(KB~�嶶tJ?�ә�t}�6/;ėO%�N�n�;3QnW/��v�ovg����v���" 7HR�o|�>�/��!�w��:xJ��@j�w}í�D=\��ǣu� �\O���S�ª��~V>8�|@qv
������ǫ��K������uOb�҅�[�DVa���b�|]]�Xa��o�ܙ����Q�(�nF�������j����ʖ�����Rf�W�w��!LQ��{���p������Ɛq�\'C,��'�%&t�O#t%�5|�5E��c�nOIJ��0Y0~������X��*�v2C�~��Em��R�����*(���{�ɟ�>k��_g�9�9�������	��r�Ws�2'�#}��>����ц���6�?v�#���/z&���^�-}ɖhG���2M�E�?>=�i�J�[W~���'<�#��˥D�mP�
r����8.�4�Q���a�~ı�S�WZm���J���D�:�D�M�lh�`���Vl�.��O�4꣐5�^2����lU�d�ة�kmr�^�o�Y�DĢ���}`�Y�H��B���ȝO�CFG�*�����5mg�S��DOn�C�Z|s���a$�f1��]�q3YL��?�������<����.qԚ�*��Ф<R����������u�ʹ��>5m>E4�������@~��QO�v���GJ�	�.뮕Q̾����}s`!�Đ��[s�q�w���G����>9��C��W���	�j^~�g�ړF�cyF-lf�������NV	�pтL�V��Xzl&�Ջ\�~���c&Ǽ�~A��:�|i�HZ[&�t��GN�"N���������ޏ���J�<��<����u���)l�"D�5@+,$e�^~̖NH�9 ��O_.�]�g��
T�����]��(���+���"��#��7���O��q�z�*���!��+��S�jM�I؄�`$�i��a��R����G/eGk�9-`����	$��m��II���J%��?f,�n6i��⇄��@KY����ٛv�����.y?�$+\�}Zlj DR�o{�%�PF[`Qc�ZZRd�z��+�Ą����.|r���z���\��ߡnpGWT?�]R�N����o�+��Ƈ�щ_�$�E�ܸ(�X,�'�;�qe.ļc�>2?r}�����l�������FO�J��ugLG�����*g&�L�@�݁��ر;[��X1�*�VVVV�^�)J�l3�ѻ ����kN�0h $;�$$\6vs�zg������O��!F�3�Ӭ�O7�Z4F�h��qݝ|�I�I�fj�9G�q�]�DGZ
X���Y�M��,��J;#`�:��m-���v��e��_���S)�H��JM����.��m|�۟=͞/��$55_-_0��ŧ@�R����ؾ���J�y9�i��_/���o.J����m�'��y��#3ԅ�ø���s|��VԂ�r���g)1�4�]����SY��7�b_4밐�6H_��&����%��] �V��V������92?���\��188A�����sR��+w~�`��2��5f�|ꟿo��=�]@���tu1��s�{�����R�й���V�#0id�O���n�_Υ���޳��e�j�i��Z�7��IE�/�k�b�R�G�|�ܕx������Hr�w6�y��t�Xnt��ŕ����f��J((�f������`��K^w�_��;H.��2�lU�\xp���e��w���|wa ����6x_�Q�ݦv�ID|C��	K���L{F�9��s����E64�c�3�ˋ�@�]	������ �q���u�'y�\t���5�7��L����G&RZ��A
��;��ն���KPp�4�z|g�'�5��(��i������_��ɭ�,v�M�E�(�3ʤ�~<�����8��1����fͨ	[��8�b��ձ[�z�%��|�v�9��A�$����e����=z�G��5Z��^��FG"���9�A-+w��l*W;�J튅��,K}K�Ą���vID�B]��'&)τ5,�@��p�����by~�qy�Q7�dsz����za˅��q�DM0 ;c���)b�1u7�v��񣈗�e�o ����uұ$K��-�������":_���n-2|;�Ԅ�>�悗�N��*��T��EĲ�傱i�e��Fb\#޽7�h����h^�$�0����%�<��5���3�(c��y�(�K�՜c����*`�1�8�6B��NS}����G�+�ͽ�]��b���B��q�l��y��{��u����W�g�Ս<�`�9�3O�`$.����v�=q�������f�F��hP��j�����"��g/綇�xP��Ÿ1i
-$}��U~2�W����sj��t҂�����^�8���O�kU�Y�F3������ٻ#�4�li$!`*N����]2�.�7�%�̐��$���j2���g���q?d��_��?Z�d���F�щ�߷6�����g�N���Q�]��_   ��v��m���<��!k�G��1W��H�UO?��(������\�`yآH�9��2և֨k�V��X��ΫVu�W<v^��[4[�������I�.=;9A����S��䙜�7��#Ѡ�X6N^�]��S!���ħ��ǭK��}߼�O��;�x����������?�P��ݔ W�cb�,IL��I��"	�{�o��K�غ�״��ך�����ȃ ���z���ة�]�ڳ"n�%��5��AW����ZՉon/�DnM=G=��_�KJ5k7�%�#荧��������h�}��-ټ7�����z߰����B�l�Dֆ�k��C�q���3mOA���,�K�A�c��/�8�y{�ѩ$���clЃ�r�� �^��i9r�.m)?�8�4%��;��h8�J
{m`}������zKla��x���m��ot���ii=I3j�⬢?��}�ÙH�O�\�]�b�d"�-��O[�C���q�>���í~���n���i�U'��"<.��V�\y������ǧ܋�zm[�1��S�;/b>S�("���_�-q��\�|�c�{�F����٩$�S�\��5�*~�U=~�}�y�NeY�2�[��X��Y��3��r���	����=�v�M�\��Z�}Oj�7��nn��9��,j8@��@�"!��>_o|�	�n��["���|�N�^7Z�Rz�E�2[yY:�]4�H���t1���˛\׍�_�
��5��KdH=�?�k}�{I�#[�W�|k�:�!'�~,�[K�ː������-�ʰ�v����4�E5�C�G�$zJ��1����I�mۏ7}K.!h�?���/cv	�J�@]�y�R��g�ľ�}ңq��Q}|M2<$obi�Aց鏵CçU�
�>E�ѷ0n&�G	hC����ǣ#V����%�A�A�{T���zϱ{�B���@r���?N��:�v7�UMjOƧ�Ri8$ܞ��q�N,�@�򹝅�������^���ڗ?�XUnP̢����IW���.��~�c���]�N�t��J�o����Q�����x �X��??�&�۱�۔K�R����+��ơ8��;g8.�g��B�O����z��1Z�;:V�x����j3�������,v��⨺�3��+���T��������~�ЧMa�H�-�������!+�P�A?� O�D`*4�f>Ψg-�� Q%��R�����)�`�H΋�hb��n��<� ++�{�,���6D0�R��j�N.��GH��[���_�sF�5�G����N�bN>�w�[�=�b���NYz�&9q���V�p{;ҋ}]#��BT%0(]�\Rh� ���:�f�M(��j�����}��Ixȶ��0��}'ws��#�1���=�\�)E��L�a-��n�|�[%� �8A
�H��F��)��V�����Y[e[������<3B	�!���a�ψW���|�]hh��͡sR�%�he���P��֡K���D1!��3/��d��ܤ�S����5������ޱ� ��R(q|��kjl `g8R��mq]�m'�����\�po���؟��ʅ��ߘ}�|�H
�;>A�n�W���fR����TP�z׃��_OQ�W���+-�x4.N��W�ߏ�M�?���I#��R����=���88���^f�P,�\�>��F��� �6��%�)W��Y���B�Ϲx�<	������nԠ^�Ԃ���PÄ.z�N&%��(f����v��r�_�y�x�N�RdP��-�&���1o�90�dTFB�c��(�_���0JXY)�b8��5�6��(O�9O/�H�3��t����A�R{zt����X'>w=D����ɵ_����*Zh�#���#y�(� ���Z�AA�)��x��0��i�O�4�#�g�y��~��d������׫>Ϟ��$r"YK����zvOX�a��>�r�0��� ��C�	�6-e�,�y���\�s���"M&� �/�x�!�R������?l���|�nN�ݍ&K65���xD�#ux�3�Q�Y0FJR�`�PSߢ�$p�\l^r��vl�T�����,��3�����WDi�H�7~%(��5jo8X�h+�Ӻ�������
V�U��D��!��� �H�P���F��%ޢN��N�Ҷ�g_��V��<KP]�Zj����0/�6��dL ����"t�Q�yF�dy���ѯ8YW��M�ҕ׺>�*����+��Q"�a�&>G�����v�)��?~B{eOW?>�'~uE# ��m�%NN�����k'8xL�5a	��cy�PUD� 0���A��ui���`�Kb\����k�?w�PP���&Mk9�l��"��\5M]�6�տ�B%�4,�����$Imow-	s���}$��;!��ʄrT"[�vz��w�g���ixy5�-K�$�d��9���/P�9h�.�x<E����,�$"EV�F�1߯Q׃�?nߥ�#�[p��	��*���Ⳑ�}�K�~:x��t�ȹ����^Qk���]BU9%ھ%�V!��C��P"��`R{����E��޼Y������$X�:/}ˇѶ)[r9�������a��Z+���S��wy�M�s�ҽ��[������5��5\�ϭy�_�QE��z4=�﷑J��M���k�d�2���\�0(uBK� "0_�"�:�z*��W&�MIa�j�r)�D�K�$��Q�O��A���-�-x�W�Fa����Bj9уi�Ts՗��@e���M֞�t��aˇ�A �����Y�;,�j��IO��#�U]�vz)�n������Ǌ56�t$��f������X:�X���p�IVp����^0��J�#�0�������a2�9lĐy�>XD�̂M�K���[D�j8�JmI����dΌJɑ�fj�G�#�/������'Ǧ��c�8���Dr���͝���s�h:՚�t@�c�r�.I3��U�ˬ��f��8p)�����i4
󤥥�"3�Z���i�{�'l;>2��K�2����m]����/E̝E�t�FTW�4�]�Q�D�ᏽ0a��3� +1b�8�:>ƽ�v��>��DVr�E��ME@zva��O+8���pp���!�^N�wޛ�w��3#� �tp�F���<!�Nա2[�2�,�'�F�ye��>����.[�M�S�C��%���Z� �Ƽup�ꦽV�4�ܒ�Ų�Q�ic���D((e�v%�7\2Ģa�,�3���S@�j���u�x�������',������
`t:ɺ�E:�gP�!Տ���xF�Ly�H�6��lP����G���U
�E����QZq�]r�H��H�H����[5Y9M�觨��FF��R��E������k.���1,t�=��S��;X�<��3��:��lP�P�53�?�;�����3�x>y�p/f(�+t2l��k��b5ʵ��۩��n'�ۤ���2u6�,�A��U��KX A��	�?������V���s�O�����mQ?\���/7B��̣Nϼ�q�d��Q�0�/7E��	�\�Ts7w�����6�tm�l�z�HZ��f�gnV%���*��~! ��� �J�R�.n5��Ʋ ��|yp.�C��/�)&$T��i�� ��~�%�?"�������G��1��?��:�R	�҉&���S�n�>a<�+�a�N�{���I�n'&^.����n���E���M�~��z��5)N�}�^�Xb������dquvȹ *<� ��~°� zfG9ɯ�j�v7�_�`��9�4�;}R��?dH�c�xƐU76
��	������]7h�&}�.��M�h�}
��e��i���ߴH�a܎�����"�w�Mk���M�7$�y��u�㶗H2@Xt�k�D��O�U���n�2�P�q�}4�E��I�!����5�\�tS��OԴ�z�r4)_�!Fɴ��t��T�,.:�vl��+ԍ7�B���X��f���$�� �,Fd���ͭ�q�|\<����()i��m��/��2�g3أm^�\�B��^����>�i�'����e���0 )��Տ&@�j�ܺI����`G�����7�Ԟl1�$P�����Sh03X�Z8ך ��j�x�S�A�2��<�WILRTFX%~ȥ�7=��s�BT�Ha���1�"�̂�>.��EV����ǵ�An��|)S�E��kX
$%�X�*z�R6_��C�ch�q��9�\��]����_�hz��ϲ�K�51���5R��ݼBⅢB�\}B�m'S�O`Θ��-2v0��8�=X�-p&=��]K?X5Xm'�3(���4��i2��3�x��0��rj�nZx3��]"��oQQS��n�Tzh�y����
h��\\�yO^����3����P;We�7�>�IZ���#k�����@.��K��iͪ�	I@��fK�oM�_���}���ڮy�͌r{�<b=rpCP�,[�٦�F3C��X�"��LR��j�E���R]�TĪ�C�C=p�l���[�=ec�R�;�E�����0���u�<�mM�V������2��E�R3*o��#�a����չ7��M�DB�Z���X�/�q��Nx*�I׾ЄFk��0q��c�cr����A7-	jg�Xm g"���y�jDuM��9��О����-6�/�{.�"�m��<�_��$b��!���uuv������)��a�P�YZ�Zq�m�8��P��y-��"T�#q��M�I�D����.�k���<0��~P#��kai��7.��v�$b,T���2�fԽB�V-��?�����>���(�0�2	�G1B�gm��j��X����P"Yə#NL���Q�y((�m�{ݏ��VWO����Hf]���>�Z��:��S�GL�H��:2��	"��ab���m{��aM�_ߐ�yg����W���D�p���	��Az��V5.?F�jO�2�PY(U-r�頩��ܧ����R�ld��e*U��OA�(���Dw!?�?S;#�\��K3�_�|?��/H5���3�4~Y�>As+P���jR�&�(5��+�,�w�=�Ph쥌�Gk��(_߃��-/�!L鄯~�ʽ຺��DѾ95�A�j�0���Mfɵ[By�����[߉��\v(��O~��GR�}/�Hך���|�f�����v�Rxð�*���0ivT&��"�s������]g֩Z
�b�JvR��O��w_t���1xіifylQK�&��a��'�Ϙ�/ux~B��fTR!��aJ�F)�b��i��̟���@e�\�|��]Ol}��7�u���h,2Y ��'*]F!�e!S�o�P)!�;4ic�7k�yNOP<�@��|�3��.��h�-���C�7
M�׹'�<����k���J�Y��A7A>����%(Zp�����s���w�����a�Z�+�W�y
���,�$ z##$KJ���@z'�P��%���Uw�V������k����$s�J2P�d��f�Q�Qd�덗XeL��`��L'C��?�I�����][!��%�5-�����u�"X�FG�(DaMĲ' g�]�n~8���Su�R���y����搥;�I����6�U���EO�l���X��-�������%�4j+p}|:I���ւ��]��z��:8$�=�I'b=@�J�%	!?i�<��5c�tp��s4��9�xT�,R�M��Fv���3Ōb.z���U<Z�����y�&���"��w.UR�Q|�g������;�~�qJ]˧XJDJ�����8aaoqq(391��P}�����m�F���=� ���҈���¯K�k�[�Y���WV]f��#���4��d�L�,�p�&��쑞�Ĕ���P�����]tP�[�E$`���2h�5�k��4��DP�ʮT��FɌBH����/�o:ߺ*/ܮ}{`74=8:�3��$�$�T�SS)�nfB-��*�S׮� a���{|A���B��%#=�N���U�]�K���!�t�����9l@1���+��mh*sm�S����L���g��-�3���"?��pu���l�G{_n*�V���ev�^.6dX�/�~�0��i�r�}��U���P��Zg���?�o�/���?��k ���|RffVVYW��*��U��V����<���Z�n�H��)Q�C��uJ��^�D����F��94H��Sdh�_�����A�G6�����dF���#z����J$�4q?; VIg���=�X:*��l�'�&]3~9�&�hӔد�
�r�}ˉ���˯�j�IS��F��;�Q���en�0j�0���nEb�ju}�5��)o�g\S�"�dy�՚��������F,�y�^a���	D�/�����(�R��t%/���Վ�O�.�ޜ,g�̀���_����}�~�],awZ 8a_1�y��Ckh�U�Dn�5�h�N��C�
0/{<f;3������.0��9�S6Ο�Ux���#ܙ��vc�FD���j��Fh,�E��T���o2`-.'FtBs[�t�,IJ�g6��*]�Gjk�� (^��Ҿ�9�[�.�����p=�rI�y�X�v��������z�
�}݋Xn$��#��5~a���fx�>�PD�b�l�M�"�,�IU�.�ej2��bu�0�2q�x���fe?K*�{����p>8&N2��ۚ�m��7��s٤>�'D��m�ÚG�|���t�����g���8�2��ξ�t�;�U�1j�5�V#��|�ξ�u_3Ё��:�@������:e����K�۪~M�	U�*0�/;������rP6���e�U����v�e�����}�R m<o����ǭ���q��A��֟(A��)�h�"!u~����yD~�a��1U����4��k��;�1'���Q$�,��^�M�a�Kn�=��P<��7��ǃ����W�ra�=���ր��A�k[;,��f��o~�������	I����ݢ7濚꾣����7������c�gBA�1��L���߾Gj�R@!����WR����0��_������;��^�<5�>���I��P�VXs%Ҕ�"��x2�L����x�B�:����wr���3�H��u��$s=�4���ap��W��n���ϱ}�*VJЀ�V����ɇ�Lq�丯���/������}a��̢��D��'�Ro�->��%�A�'s����,p�]y�Ft��R��f��������=q������Q3���b�9�9�p,-�E�Ui�o�ȅ��7���=�cT�`>��G+��P,_C�f���/�9v���lf�:�祡��p� ���iDx�ēN�V��_�P;��ݡ��z��kPb�g�'�.�m2:�F���[j�F�?�pe܁�I�� ��[H����b!5�O-,9��Z%Qd�)���d���O�Q��0���h��O[Ø��q!�IjM��k88���\j���,���}�T�p�J->�Ԡ�%P��$+���V;럄p)�!M�����H�gX����F��t;���H���m��U��X�¼�:��`8����9�H�����`�Z�rьf.�,ޱ�x��LZ��ﱾE���f��*�7����Svr^�K�3�c��3����`���E�v�rg�rf�k�]�2��6�<�jG���*�l�i�lH�F	q��d�E���Kp)'d6��U��5��[U�zKRu���zo>���>�ID��y��{`� +V5V2"KnG� !�����ld����(�Y���yZ�����6wZ��c�h�v�c���a__�=�Ѣ����k�`|���X��m�,M�}.�B!�D�Y�Ga։���zߤ�Xm�6��X��۝O�h���q���Qw@��(����=ߡ�$�"�����q��Â@�a����� �QE�k(-��h�~��DL���	�rD��  �'.fw���`��6�����N"�Vh���s�@cV��s���1����S{}�/��'ꞓ�$Ьh�5�"�C��v�߿���O�@��lO:��ݍg�8�rꝗ4�Q*
_���W�v܄��ϟ��	�|=X#�4B
�6�И`5C�XK`X�c{4M��W��8˼�a�G?��b��K�¬K��6(������8�����/(Y��ݏ.�Wm�"�Hf�e&�!�ϫ1-���xΖ?����pj���SX�cx2�{�ns ��%�@V��%T"樬L�._��e��e¡#�G4@V%,�����n��|�:�H)b4F�������m��V�J�<-�ҕwPF��M�I�1�?9;�DA�����7:�vH[�F� �<�.6�M�B���� �-���n�ʬaX�Oqc]����>�R*��'�����z��Y�wU�S�Ad���q	PXP�R�i먨��K��)1�!���\\ބ��� v4L=�o����:���_�8 c�T[m�j%�%��?���ח�����T��Ge��pe�J��iu��(�" u�ݚQ����!&�'�����q�ӥ����Nm��b��Z��`uyRuh~_{,��c��d6\��2"�\҃�e���bOeqI�p�8J<�deT�fշ�$(�?�-�Ջ����ǂ����J��2�YӰ�ޛ�DfMHH����F#�\݃÷��4�ѡ �{�W�*���-���0z�MPP.�m�pbj�m��4X-�a\J������4Ͻg� �����&�$���H���/`Q�ʧ�r/��Rr�~�82̒�E�����؋#����o=ߝ�'Hg=���~LI��cF11��M�����RV�;���pc���&�^*�f�#W�Q4"���!ۍEƉ�>WT\�M����M����ړ���J>���Ri�K]���
�*)�W�M�3/���:D�8PC�f��5fU�E��5	�
��)ľ��lN.�>m햌��QCrYJ�B4@
�����(ī�����3d�AD�^n-���eg-���d�W�(̢8YB��"�N�+*����Af�oh�*Z�s0d	���;�۩������֌G�v��QT�M�Iɒt����3!���SW�Zj�WWZ�;��yj\�&t�_B�6���U e���kw��!e�Q��h1��N�ط��eH�O� 8��B�/ؒ'�^��k�*��ZgPc/�\�˃���*6O��",���B���0�&�NQ�88�a*�H������H���lRh�mܚ�H� P��1p)�IQ󯜌g�S�� u�<����c�c:ݝ�����Y�:��*6�4���W橛�&5N�b��k#C}ߕ5��� ��o8W���;���ۤ9��玞�[}��h�Ŵ^�lI���R`<�q�Լ�� �n&H�!KN����Q7+?��j�"� <�i�y��2\�_�ZZ��i�T
��G�5)���cS�jp���Bt��|��T� ����f`l�f�˥����_c�KL�ի�xVH��:Q�8����橐i��L*�Lۯk�����/Q2���f~�������q��zsw��g�N:Ae�_z�Z�^G��?�-�=7��9�����]�MUB�'�I�¦����Lr'}��=_���_�����w��y|MW����{3l/���i]��{,���*���dV���?���x� y��k�����}�E�8L�vի�b���?��˙�5�?-����C:d~s0����u�Ӻ�'��4�FiS�-�$䕋�^r���,���{�=�B��a>q���p�o'y�,.ʱf�r��P���d����~�@-�-N�kW�6ό��K#�Xk>U��<Ѐ�&�%� �2ʏ���ަ���_|+�}���z�ҽp(Xb�'�����G!�|���4Ku�t��4$0��c{���p�K?<�m�T8�8���JO��K��=/K]��冢;�=�ڿ����<�=�=�,x_c���'�yg�W��IvT��� �;�`�����c�`Y F��n��-��xû+}�x�O"�5{	��S���e��_̑�ԩ�qhմ7�<����G<�?dػ������D��g=¤��u�do$Uv�](�$Ϻ �-6�F�;2�֭��3SʲT���4��D�c>��*��)?���p�� �տ�(�1�0�����#�Ph2�ed[�� )�����L%~N�l)�!J0񹄓��qM��'O�<�L	�}s�m�Τ�R!IzdQX!�����.���	��+J�v���0?�EZ
��17�k��w�4[�<A��b�ߟ�(�~���4�b�m V��V�PdRW.+/A���Dq]���Ԯ�w�ۦ��3�{���}�HʔM������"
;*A����wgWte*�w��Q�3��� ��ޞ�I�l�\Ѻ�0�2�c�b��N���|�:E���_VG�	�\��MǨ���uGJ�Q$�Yy��_3��za�.�tJ�u�)ױK�~����:��!;~5��䟸{���q���?f�s���9Sx�r��6�^M��Py����G@7/��P��=�*87���RW�����Oz�sQ�*���,�4������`�����!'S�x�}��Z��n��U/���'/<��d򯯩j�	C��(�������S.�Fg�y�+��b=VHkM{U��[��[���v,�5M���( �}�HBG�,��*�Oؒ���ڤg��6��
9�׻3�k㒡�q�dc�������1"(�z/���-VH���Y1~�J���kD);�񩩛�~�F�]�bu�8
�kM�!3��r�p2du��5�4`.=��i98 	m�-/���0�zf��}C�3�ɋ����@��g&��4�6���H,��dկA�]`zZ ASK+�9�]�'�3ܻ?sw\J�r׮�)�'�W#����_��53�d��S��� C�h����>�=ƬL&��^U�c��+�8��[�]��j޽EǸ���s/�{�XX��A�ɲE�t���R���s�eV*�2#ƬFlE�d�o�\��r7�(ǹ��|^�D���&��n.�w�M�Yc&��i�(v��Pa�������O���dR$��ؿ�BY�ѫ�#�j4M��q��š�%�"�O�MX=���mNSb�Y�5H����)aA��Y���������Z-/�(GK��N$SG�䙢�|)j���5�����[w<r����b�I;K4�6�+�v$����i$I�e����?E16y3y��s�ȷ9���&MdG@�E!���2��A3�!��̡bP���dlx�Q��b����R�x�h�b���)9��.l����}3`��_�����(���R�g}�M��2������$c� M�:ݐ��4a�o ��k�va��@��C���)�f�X�]��T�[%�`&��-M�Q)q����M:�F��{C)���: ��F$f��bkT]�ʠSRS���������Abe2�}o֧���+,��*=�*%���g�Ͱ㲒�(oX��j��;��Tq}K��fE�mE\�(m"Jڱq�r:�=��sq���t�o��,M�|Q�U�8j��le�J��Ʊ��к��y
U���BL��fGe���/)��mEN>�.�;�O�uL1&o��Hߥ�kÒ�R�S�r������ ���1L���gn3K���XT�򱠒f'������X6�y�}߄��v���h0İ5�7P��Q4@|���k^����GJ�(�w�ڑ�uZ^��)+����n��2�D*W5���',֣������w��`�$�����X���ʁ�����"Y)zCa�LfB�>��F 1
* �1�d� �:5�53fH��}���){$��DԔ	�q�`CQA�<�֯�/O����Ϟy��9��jX���J��,e�2�(,_�:=|��.b��<~����~kH22�ֽ���b�1â5��pg�7`S�hD f�|��9�x�mk��JE4u�E�w��綥.u$C�� �RLn�PN0Ţ2��AL�|*+!�]�SX%�k����V>Ysy��"�j��L�%SoT�NɉT�
�ź�K��[��o�e�^f��H��fF[*P0+�i���s1�������N邝յ�/Be� �ǰ�0U��RUWW����� �bѐhXE�hny{�����!�Z�|��'��4=J
��h�`�cՎ�Js�T������'����?���'_L�̲qSdK~E8ͭy.�vt+[��J``Ȳ�Fq
d�t2��v��3 �C��n敟�z��lU]�g�4���8K1��@&�r�$��n�;�U_�;�:�ű#0d0_��,w��e�e��<_m�'N"��,v��!?G��xG�n�
O�7��?��;�%W��X�0��zr2 �|6�'M�"�O�hP��*�̃SH1��^+�A�o��;L��=a�_:uJY�,ƕ∵f��/4�}���o�I�:N��R��G?���Ȉ�f����
R�a�R�������Ĉ�m�ZA �e���6QRH���.�Rc���фH6��g�5N�J v�aZ�b�	���\����E���[�"�6"
�R�2(��V%��[Pl��l}+���E�'�.�� aJnw��"�Dl�(����E���X���[^vt�}��f�R��+@��]��3�����g��t�W ���o�$�j Wo�V��F��˃�'e�=���Ȅ�d%K�Y�vh�����~��8��D�=�ov8kv���@�^W�<�_��V殘+V�t�bX�Q�Tu��[/&�e����.7�'�h�@��' ��K��K	�ř������h��	�۱�:&`�*��2��5C��,{6�	�T��tW�?>��~{���'�J���c�H:⧺�V���gcC�X�s^����A?��z�=%� �B�\I�lJ����!C���B��n�P�Y�����r��lhԔ������Q�)�v)�K�͖ �� �m��x�m� C)��a��3Rd����OMs'v�_}�<�����s՗�#p"2���[\�)�,px��I�>��XL�$��ME4lE���˂�������Ɋ4S��[x�>��6_��^��~���4�#�/�x��*8M7�@�XKʇp��<Ē���}���-�l�(�2����4�y�=Ę�̰�{d�������\ɀ�7ilHH���?'O\���G���R��a���Y�L(�L�V�~K[�T��<��I�a���~�<r7�8 \J�:e��d7P��EF�%�n�[0���n���:Z�>��o4��_Rޟ`�!�F��y�i�W����t0$�Z�F%�ygu�O��j���B�O�gJ�%Z�XS �xe�k�ӘH�
� \1��)?�[���	��z�����I��#�NbD//j�r����/ז�i��Ƕ-���A׿J�8����w`���u�c�vұm�ݱ��ض펝t:vV�۶m'��sη�Ox�cָk���	��q*�QӜ�B�6�M�c�Xy#�-��ݫ�J3�����;}M�W�DQ��,�D�}B��3�P�x����X���G��b����.6�Z_3I;S�;�R� #RS*��Z݉W���(�y���2E��7`>������6k��3Qk�D[�t�1U6T�.��ܯn�����ϛ^��͔�q�R���ӈ8N�v�ˋ'����:��e5"D%�}5~�H��j������rc��}c�ƞp����4Y�:Ur��S�/ +\P�o�O�D�h��1%����B1���)�f'������n���G��O���!���wK/D��7��_�x>ݡ�	�����g!4�y�lL�G�'lǀ4��2�
����8�����{�S��a�L��X�������ǚO�C,��;�ے�����XI��9Q��0E(���&B!��m������ oT��� �`0P�J
Ť\~�:2��˯�J��FTt�l�sE5��ĉ��8gN9v����G90B���y�N��\�?OЈ���
���x`��թ�H.��h��y��g�%���R�F��$��-������u���多�7h_���U�D�>��_���2�mF�k���ᰂ|�B܊�% 赔(&/f�b9��-!�}e���|�z��j�:�Nfƶ�l�6[�>�NUH+���O���9JQ�$pB���HCi&#(����Q���I�f���<�v���� �ZJ>����x��b(���^q��1T&g��K�H���qBmn��I��~�~��h�ߜv��D\�W�wce^1�A�Ĝ��ԓ��ڐi+-��e ��U˘_��0n�.Kt/L�yn�lM���i�F�[@3�rq�3��1��$VX��9ưG�ʺ~��"�D�˺ăVp��99
62b�A��}Tq� v��fch���V��d�/�\D�Ӥ�m�	�/�&7�4~w�0u;G�ek�C���;��O�%���g�<��N�����}T%�n�I}��k���t�cҦ��N3F�K�ce*#ooFic�A�� g4�a�R5Q��(�wZ�+����S@�����Ȍg���<z��^!�����Ζ9�����{X��4 ՓT����*}�kFȴ?��}�Lh�8#�9�D��:z.�x*��.:]�!F�(�����߻J��y�=�\�W�w�~���=���|��lT�w8�i��F�A(�"6~�.��b����_|�H!��?��y������<��wʝcy>�{�r������a8QP9�ɦ���o�	�uZ�������WGC�4�oI�
�cYZ%�&�!H[�G���@G�҇w�#o�o]|�ԓ�[�O���Z6Fx:�����	�DS8T��ҕ�"��>��0U�m
;��ѿY��g���ƘF�C'
��W�Mr6�gm� R<eU+eiԡ��e(�ۆtn�k�ϵ�wbf�#�欂�(\�	��?It�,�T1�!�1�GLz2	b���<��J���td3�@�jq &�1���$ݒD{�*�g�nSz�z3�!�?���{��T��`�@�M�P�:�2����;�Q(Z��X��g�F~rFGJ��D��bʚd�#e�,=�[|�}�/��FR�2������2QFj����;����!q54���ҕ�^e�tɏU�E��@B���>7�:l�0R�j�lST2
L�E�w��v���$VD����̏5�'ަ�M���f����Y����X1.#i�CD^L`���7D{K}α7�Z56M��7���vӟ&�����2��?�l�v�({Y*L9��T?s�
�~���_O=_�9�#f17����e�鈮�d�NG��K�񛫟1�Nf�,8J+�PբY���O�� �ѫ�D�#Q��ٲEٸV����g&,<X�I�F��tj���.�3.�+G\|�`�١t�uIo�����*�>���$���Ae�@��1^�<���
���v�ƠC��#�����:��'|	���nFJG
4�xK��QL�Z)�=7[{�K�f��(�2�$R�̼�)~����됉��U�1]��3D�+Q�n,���7YI`(���r^4D���cbY��	/�q};���~ơK�a�u��=���{n��y�����`�d���_73kP:ԩ�U��Q�@�(PѭOn�H�� �xS.8����y���f1E�7q�w5��s��hK&��f@A�o��(κ������z�I��~��u
F7�jPc��qP`B��!i�Y-�@t��*�����N�z�:8��?��{����`�ڰ,�ʿ�2�aS0��k#gD��ٖ5@u�[����ՙ����q��Xؙ#J(D��	u�{��yyrL�U�|܃������×���mp�:��h��ɻ����'�����8�L�ͬtJ�Su;\��6�߾+�O�*��[h�d���3܇%�D��XƁR2y�m�U+�P�����+�����Wz�L� XUDH<���!�ƑE?�_:��y`?��۲x,(�$FI�F�j=�("_�(UR?~ �f�ʸ �8�4rǎO�a]AU�I��Ԩ����Ƿ��Tl�L�G�Ā��f��o��+!�B)f�t��7��bOc2��z�!~�q�$�RW�0Ӡ���ƍ�b��2O#ĤhUz�<ݔ=}^�����Y�H[�:q���`^&iT�l�vW\Y5QwykV��'�iTT�O����\4��ڸ�_�8�,�"!7��X0J�&��,�6*>"�Ȉ�j�l������n�>+��V�Q-k��ي��$\qj���Ϗ�
�]N� 2�5y�%h�  �^��Ze�y�u��g��]u�Y�V,^�^�E�k����v��\���_1��X6�����4��N�=:|�x�6�U:e*�Z�?��}�z���m�؜3�����9�^�鶧���]����>$ͱ�BELm]0����O���lW��.}�t�*�(ߏl���>O�U����oi6l-�N9%�x�LwECy�f�H�(�\��oY-�V�,Bޡ��a�B/j!&l�V�n��d}iT0�A$��KS�%�p�{�O#o8k�|e�נ,�VV�p�5G�G���N�@b��]f��OV-h�|�#o�<�+&��x�N ����d�`���?B,�����;U{4�CsHՖ=�*���0omB��6��L�8+�
�|P�h�<L�.�dH�ҲuAõJx��x0��rz�Q2���pS�@Aѕ���]�ftH�t�Ϥ���N,VJp%촴��<���じXf~N��b��:f��7��Z0eNm�'+ ���2Q<� ��SQ��O��3��	H�x��-��$%u���|ד�&}+=`d�#�˵I�ET9���)���`��;�|�,��=l/�j��4�������]����@Q*���@�4b�O�)�;���e��DE:JIn(�Wu��";���7lm_���?Ɏ0ڮ�̓=�B^�C��z��B�:K�s�
�N�ώ�/�����z�'�Y�t�#��4r����Ȏz�&��挵_�B���n�#� ��Fq�`409YQ_�?]��'�t�Z�8{�}���|�tԱ.�(
�CGv�La����+
E�ڈ2B�x���.%�O~�l��?͏���z��P�*l؀\�mIv~���V�/�5����=��ܜF����.Uqq�c��Y7쏲�䩣/[-��y'=��g�>TBcx/6�Ok��'Z���i�U��IV��J����y@T���9�23������Yv�Ԩ;�l�o�r���݇&�,+\����<�1J`MD���n�[�&��W�����Y�������j[[ǹ�_�}^��sFN����Ǆ��G�Z���b���Wp���|g���&+r��K&&O�a���Ɩ��eVW��G��|�$�$9�\�
X�q%��vML>bDׂc�<��ޑ"PT�i��> ��8G�٥B�+�bv[cX��ғ�����+eM���Y��
�@�e�����0%�ڧv�/�;[npG~���Y(�%�	Dyrk����P�^.���cf��}?�����1�Ԛ����y�薀�-�N��K�1���JR���U�;�Z۲&���2_���|��G*��z���z�sI�-�LB{����h��{$�	�h�CHÔ��$������v�5��Qs��L��ЂLX�]�Z��s;���Bhl{��ub>�(B5�e�'9��7X��|Ĭ�#W�3�t�C�_?1zQ"�3+�xW5;�"���M	��uM2S$���9�0g̥>2_�B?�7!7��������1X�q {�;M&��KY�cIR���FJ�P�ѳQ+��	<J��Z;c����~�m�!8�x쓉��.�cuX�c���w8���ڸB�bINN޿R$���Q�T��j��213��w:�842N>O�Y�EE�|�ñ��MS�q\'��6���8u�PXh�A������1fM�'_kD�1�뫯~w���eCK/��^x��	�����
��%(��e��/G�]
k�Qb�9�i��ѳ�3�4d!��ܐ�B#`��6�H��2��x�|}����w�Y\(����v�\�]+g�4'���QNL2�Dr�˴0��\P?˹Ռ�4�'P%8��e��!l�U���Xo�5)*��@j�h]�K����r��OV���luyAs_w�6�8ՠyHM��ſ�~%��wN�?G�ˈ�{�[�
�b�?�a+!$�H��Ցd���D����kb��?nU��]B�|�b�^&� 2�8�e7�y%{�|+ajx(ͪ+/BxO�ZȫwR���Q{C���z쐲��SL�7��>�c�ƿ���Yj{T�p����J��T�g�zlT��(YCY7GY-i�o{ʈ���:;nG�����g����j�Q��u������x�w��+��7�*����	�����|����#�-!+2)���U����S ���i�cY*
��k��.C����G���˰�ʛ��i��������H��%�U/�r�CT9����}�t�Z"�h�������������qѴt|uU�I?����d\'�2���
���#�o/a��. ���hbc�m^TWP�ڼ0~f�m.�p���U�fڢ���F����i�f�����W�����޿��⟛�3u�ұ�*̽�|�}�WL	ʱx_z��P4W%H�K��~��ovfi ���H�`�Z�$�_�5S���ۥ�����dQ!RJ��t�y�s��+|R��6d�+ٸهs��A��[z1qq;o~GȰ���@8 n�=� 0�Þ��vP�����ST���.5e�y%y�I��O4�$U�"�>i���Q��%����.M!mc/��r�k�Դj�>s�.���s�=t�Ut��tw��T7a���ͯ_��#��Z��
�RV�y���D��3e�e�/�T�V��}Q�C7r�t:�����b�7R��p��X�Y$�j~T�����.��4oB�����3x�-Zo�G6�ŢB�1&oe� Q�.9&��˘��	$�s�3/-�g������L��lЭڋ��#�����Uw�(v���9&=��q�e��:�M����=�L�_�.��ڍ�j�I��⻴M"j[�a���D�:�����8Y��y����p��ޕj�6����0��˳)�g %=$���<a)6m=���be�6nI�����=2֧.OL*�f֦�� ��ߺ�X�`��.8X�"W�_�x?N�ά�"elV..�6̾6��=>�����j���q��U汳�>(N@h��Gs��O��y�y�x���$�?`���M@�pנjX;��v����z�/��Bd��\ss�[��>�����+�2��QkTY�F�^��J_6�v����F~~�#p#�Ym�k'�f@��Ǜ�c�"zhJL�腞)~��
� �&\b�Q��y<����Qg(M�Z�ۺӘ���˗=�X����Y��SC�:�V��s?QI��`�#�s�E#9;���F�5#4�+����w�%$�k���V��/PǾ=��s��z�+���r�ڴ���<���u),<|�����u��[p���o$�o����h2��Lъ��Fw���Z�&�D_��%FǮ3c;;g'I$[��&#T~^��F.��*�#K�k���'ʪ+�Z��I��\��V�{+���[=V�8��'����_[r3U�jo�����V�i/|e�6��<L�2/�g\X>Y�r?z�Q�X�>uܻKj!�j�LfS�4�~�!������
@ 6G�m�֕���\�'�ʜ����병<cz�M�H�J��>$e�
S!X�/�����_&y�w�q��*:Q����_�w7��|�b�!�潬Z �Pf6�Kx��7B��{��v��{�N��y�?��Lfʺ�P �W��rU�z/���4�+�*7Cօ����<��p?7�D�5�z��mR���3����Y^��b>����j�1 QET������⌛c�R�Cq�e��������g-��/cĂb(��#�X��Y�(IS�fA���'�+�Gz�K�﫤��NE��2X�ſ/s���(o$�9���[m��^m��V���f����n�;H����<�m�M <)ĄWM�Ź?���Ҝ�8v��D��7=���g��UK�����tJ�mVꁄ������[�â��~�m��X��[�g@���v0r��T�����ĒVT8���`)��J���w4h�UqF���W��n�P7s̵�+�����#uh��F�J2`�@+)�Ȝ�r���̐�^�~�7A�\f������)�[�l���I�Q���/�?i�2,,Xn�!��! ����(�È�P���R���T���m��ZT���zw�)��_(��$���8�<ee��&%�+�$�9��5�?�	ٛ)�S*�DK�f�et��io�V�A��U��ct���y����W��[�)E啔꜏�F�G�o���?�-�+}ڲ��gc; sS
�~g�M��J8z�9
.oHQ�X���,���&�u�ա�tb�Q����;��{6���HF��V~�
�R"�54�����A�P�����=�_��F�~Y���ѹ"�y�Pk�A6�kd�l���P�Ak��K�l�ަ�T	�e����7��er>��?e���#���.c獴�O�bH9#���i����,��Ԅ�GP�ݝ'Ol["����pV}eb�s|%#ӕ���}e<7OSu�%� ���(\(�������-�:ԭP��[��@��c$d�@��.��/\�H�F������7�2ކ���dC��y�B�$M3c�V�W�2r�J,( �N��qϨŸR���"��
�y:&����\vzGQ8��������wO�Fٿŕ'`f����4���(�/�z����>L��7st�)Pi�_��f&�j�=��R����rKyY��=�=���^�S0����b�m��I�8�ͤ�Q�u�r�lv��\��
nP�	�uͭ��ƂH������o� ���B�����0%�,�T�ƻ�qI�(��tc�i6��ɿBi�o�N��[����t� ��B�˱Mklf��*}�?�s�s^P�c�d��1C��ﲊ�­�K3����'M߸S%fA�M'�0C���gz։�B+0S #�쒮�;��b�S�p�Ø���CJ
#و�KN��Ԓ��y�3~+Qs|sh�lA�T@Ն�1�h�������a�ܩ3��<X|�77������!"l*U$VNɟjuX�?�-���� ���`��r?GCY�$��ax�+�B�:��5^ݻr��E��M5t�Y)�P�����
{X�$j̴p�ǈX*�pڮ�L�/s�B��4����<c�߷�u�ȣh�RX��(�^/����?���#�E�E0�ٳ�\�K�}ł}ܻ&�c}�n��WئX��6,�qmd`��Ӥ�籏fࣷ�J�B)9��ِ6�a]ǧ�����Y�y&|��RE�c���7��ǟ�Ạߎ������sd�� ���J��~��t|7kt6e#�;�(�7��	R��$jf��/�!sJ��`p����{z������Xlm�����o}|oҎ~���|�mt�*�e��c&����-���?l}�6���\��a3����x��Ʋ�l�b}�zqY�U�'-7��c��ʅ���$*1��m��gM�A��!�Կ��ZO�|v.l���64f��80fH�����}�O�+�:%u%5*Z���l����!���0�h�럪�K[Q�%4j�(_�9����Oֽ-��7�ʆ���m8|qGRwj�1�39�����Y�벨�����<f����=l�6M9}���l�x���yZ�tPb����t4I���5������ �+'�KW�olOt�o�x��fՂ�?�=���^�2�g�[���o����f�^����a8���4Km<)��4�z�@�]$J�9�c��FӈwS��W���#����g7?P,��E6�(1�f�&n���וY,F�����������Q�f�~8�2��C��[:�q���V0V����_��b����D&����T։�ԧ�V�}��?��n�S�����ذ�YC�-�/xڜ]��_'_R�̏�6Ε�5��Ir��3}σ��^g��|C��\7�&yfm��f��B}[��<�Z�~�t~��}6�+��j�"M\o�ߏ�wL�P��ߦ]1���@�'S�H��f���]�h�h���9�%��j���8	X1��!F��6�.^.�����UJ7c5h����p��1I��>M�[�L�9ˈ��z�7�mZi���m�4�s�8���28V�5���d�8Ÿ�j)B�MABJI�A���\G�pΤBO���q���4�r�ͨ2��J�����h���lHy��ަ^���/��1�^ċ�9f
��9Xnv�kY��t�r�\��䊟���ki���k��,#!���ǨSIR�,��~G&>��tZ!���Ǳ�����|�)IS.l㔁�PiC��2��o���G+��׳�t����.r7+$Tk8e�Q9�m�'�˒�0��'��}���s�[�OFO��S�u
�k���?�r�q��x�5w⮦�-F�A0_��$?++�ĉN��3�&v�ż�c�fO�T�q���d����R=�,UOO���6�����n�3E@ON�L3���t��9_�
�u"�����R�#͛J3�!�6�=v"�AK��5�뭦�_���⩺
a�A��1��L|u��n��z�Er�[���R�w�8��M�X8����/��ԅ�qY?�����6���߷{�bA�|�$�I����u����?~��pTLFȕ��0kgh$?��EO���6α	0�EI�����,��ij�R�f��#�V���oM�eq�Zk��O������������a'�DF92�)�6�}��tq�ч2u��=3\@��9��N)�	}��@�����X�'Ic��.�b�T�i�Z�YYF(�~:7���+��������c�-� e>�� "���^�2�����z{d�d���i��_g���P��>@d%�d#���]Ze>��Y��e�S��4��?����SIQ[}v��Xҏ�G�s�_�"
q�W���=��\�a.�l
�Zu��YYxF��o.گ����s[r=#��8�*����x�o�!.�:F��6�)�.��}�tZ	9Wf���&�H��4���?�*�V��O��}֬\,W�u����RPL�[Д���k�t$04���P����Ϻ�v��٢�����ۍ�ha�5m�(���^�E��>�;1#���{F̊Q��a�����ݦ����>yHN��6g��q=��
T8+�%&�����f��O&� p�K'��|Ǌ�)Ք���?��~�A���.℩*�0���Px�d��h�N�5�:�3�(_3�X,}�MN_J	�8��x�2XGX���7g��w0���/tt������H5y���XH���5�1�^ք�ڄV���,����vfg�,X،�F<���hgo���-�y�w`d��J3� ����Ŷ�"��/=�C��Ŕ�f:X������ި\|�z"n��I?�Lf��I�Ж܆WH|H�����F
Z�=�q%��z�.�ڽ�^э@�00Ax�1+	=���ݥ�~TF���6}@�wgw���F�J�����������W���!���a�8fi�B�V�U�e*Yi@�tX�֭V�m:9��;��/5S��q�*ɑ�0n�b����l�$3IY�>������q�\C�,�-�sC�քY��	e�l�l�&����3W��?��G�cc�����]c��6U�;J �ߧR��9Qc�`P�"!%%'_��Ȑ���+
�MF����S�.*�rޞ O�������R2L�(�C{UN��N�h�j��ǫ'��Fc�ԙP�����@,�ݮ��p;l���l+!+S)��Ҭ�,[؏C� �QcM{:��q�����sO1�HT	��l4�D��w�����zJl�4���cƝ��/�\�#�7��R��!�a���R,�`Nf�L(�s��U�(�W XC��3vwC�jj?W�5���*����|O��v���1�7�ϰ�D�bIg4ؽh��=x��E���KV^ޠ�7����1ά~u�i��F�`���p-].�f8L޸��ݾsV�x�T���z�����{�vh�'��<Y�F�-��؋x��)�ZrQJ��u]�/��Q$S���e$�t��[@r��(g�S��������.<���1,�m�KL�K�_%\���5BT�x�?0m�N�D�z8ЖhĿ�B�A��%�,�+)Ɍ�i8�C
��kI���g`h��u��߱���7����:��R>M��.�sG�m߂���oڐ���˭�/icf���A408�V�xF����/"A�AG��NҔ�����3�3yM#�8���7*i�6�n�貈���',#ON��@���~�D��.ZzҌ��9z�h�֕n���f��ʅ�t2
�b���k����+�M�HY:E:�<4�� �!kt�����r�/V���[������jF?ԋ�� w�F�DKn2�h��48�k1�mT��v��g�1�\3~۟�?R஘tBL��Ԝ�P�� ��F�e�U|���)d�p�[u�4*9C�6��<t
`�520Џ��U
ZS�Z�SSK�p��}�e�#��U�a�qW��u�D�s�0F:�Uw�j����QL?|�Sá�I7F�}a���Mh*�L�:�8���SAq�`��`VLVV"s����/9l�|��!��� �rs4g>�u�q&FQ��7ĭ��w�׹gzO�D�ܳۚ�θX���ȇ&�P2���=���g��+�_fQ���g�|-=|W�{B�,�ļ!?i���i��z��g�����W��4ӂ8�eTWy����^���b�U���$���ED%�ޒJ]<���ao��S�4�?�i�=Q�t��q�";�a�� _����!�~�<IG�@\�(��g8�%�Sh==ɺ$X��k����zsi��-9,�U3��j���V�G�/�p�qY�+5h���|�Hp����7C�d5g��\��[S|N9��ܭ{ouJC�o�����N�7'��������2��P�\*�
6�[��嚟5��y1C����pY������V˺�����ob���D�U�yD�-C0d����[��e?������ 9x&����޶|�JJAK���R�	��>�/�$d O�bЄ�mS������S�>�Qd�P�������e�д$Mi�d�� �V��F��0)b_�%W-]-c�1����P5v<��h�])��08`��L��bD�b��`�Y��y�����(,��6/Xj�da	�삾�qƫj��	�<��,gxE�V0X�!�W�q�<՘���X��!��K�x	��*m�rC}}��9=𿀕�mV��pi�Mo����u�"Oq
]z�&���4��IȠ��)���M�=�Rj�&G�}|WU��G��������ʼ?lBf�=N�V�0�}���@���|+V7e�=<::�ݤ)`8���W�2�՛�!u��u�ɖ�m�j	�ӎ�����}��u/4.!��f���h����S��=[�D�'9��:x�J��
��9b͚t�"�G#CGc��" }.6ʤR�Pw����6����\�MO#s��ʷ������I����Ue*����n�;�˭]^�]��q�F�|��@��v՟j�х���0h0	$,�<G9S<�������ͧ��dl���W<y��-]M]L�
~�U�TM�=([�^n�2r�DS��>�=�w�n��.����b��U����'�6�9�U��ғ]�V`4+/�C@���w���w�N�f�"VBG�z%�h�m��<��m��\�v^�Ư�r@?}�u��w�]�j��?]�t��|��/ݎ-m�t*M��=	
ӡh��@�R�|Rӌ�?��_2�#S����n�s��z5c��`��:�������|����S�C�Jcc���I�餾rq��VM�=���]�9�||�BM9@��ddz�(MG�J�k� <���N�}�î��1��������d�����������ˍ���3S
?b�@x�����m�!��%�����)���+v���ܢN����}әB�]�}�*��Fh���7G?�v���~�S^Yt�<�*7*Ʒ6d�&{?,,�����fqȨ��G�s�ߋ�&��������7{�8�0��2��;h���O�{���ALW쭽�}X��ޡ���j�Ar�	GX�����a�~�]��O)��3{|}x��ZWʌ/&>/��w���|����~<�E�O[e'�y�x;]u��3��2,GS���_qY@ϲf�Z��20��k�*�$�;.2���sq���&��,Ԓ#,�iή�?L���8wn�qw)���ƌG9i�*���}qu󱢵/�j�PF�dn�A+������*W�H�{�y���룥��RW،��2�Z���I�=�	�'��̗K]�M�b����m�����<C��9-N��B�5Dq���(5��.,2�uN������sG�3�xP*�y(�:�V�F��%�{���o|�J�!�u�J�����P_�٭� ����h���v�����v=�h�Ԏ�T?_�ObV{a�2���#6l�	v�+[�}�+�6 8���/�(��)ݐc!�r�6���k�.��넶�tROq��( �4����:=ʛ���	2V�Ddd��>5M9sMRŵ%Uࣁ�g��M6�A%=�^#�I�z���Z�?J�F������< t|��W�<;h� ��B���AFS|P%�)�f���J	v�?7��'Һ��]þ'�������prr�F�6��N�R�q\ka����u���#}>19���ޜ��6�Rk]�3+nGM��:o�C�cI)`H  ���ƀU��o��F���\��I���b��b�(9f�5\��k��p8l��lLm.?C���Kѻ�Q
]�`���;W��1��j�j�[8��������������1,9�"�wV���8o��ݦ@Y�CiY��w�/X1�=�2�<�37���A!�M��xԆŝ�|�Y����ͣ��xf��Ȏ��F��Nk+U3;��s�<v��s7�\/m�q���G�}�>����-�a����#�5K�?PlY�y\�h��_��C�?h���r�߀�9��} [�"�H3r��C��ص��	�v2<��IO%�z�-_�/U���m���y�҈��U�h�n��S�(���3"�Z��\s��
*aG��@a�z�g�@	ح>�ʛ��,\�nn���El��Ȟt��\��PŖ@?0�h%�K�,�J�����m!���m�Ek�`�ʩ`aI�*��%��;�������3A�5�[b��Z3S�, �r�tE̱w�.0�jJ����Ĭ�$���j��%���q��~�xh�2��`��B��l:_��$*��q��ͨ�����4�[I�(���ů���þ�1��e���H���ro�Ѯ����V˦+5�� M�&9?�>� bǗ>:xs�ɣ׸����d����<NH]#��4��e%����w�?�b�$u�RՔ�i4�KKkn�ÔT����܅'�f�-9o�F`����4		8���w�A�r��*��4�ऎ��L_�5��%�/ݑ��O<�x� ����Q��\�>���]��1��<��42YV������}��i�bP��	2�m_$ԡj�E;�**M�*б��j�����>��g�Er�E�U �1%�"4�li+/Z���k�^���\��=)�ׁw��������='��o�6���#n�a���-.�vi�=\��\���"Q`U�����>ʾr�o���n�/I�LW�m�O��iJ���*Z��2��B�]�T�M�
-���R��_So��-}x�XQ�&;I0��G��`�����׷	p���_����{ �w^�g Lv�]�ʤg����;�4�H;�Z�B���<Q�"�[�]�t�vc> �n��aw����\�Ր�m�Y԰.� ���6[�*S��:3�;��ڌ��Ec��M�q�ݯV�}� 6H3:*gY�L��l���,Q_���U�$�Uւ�`��B�zz�8�$�ݵJ�b8��͉�>7�	Ʊ1��V�>
���KP�Q��6��N�����A��a���3H��M�b��WoԂ� �Z1=�p(t�*wc���sX\*��1�T�5��O�u�$NؾV�;�\�B���?�Yz�t�+䚊f���/`�5���E���+����.�/�0�h�8ؤCϨ_<��g(F�dP6u����Ԡb���h�gR��T~��c�Y���uFf2נ�B���,}�p+����M��ת�Yq����c��w߄�����X���Y�J�uJ�=PO�D�*���`����ɪD�3
p�B��eC|���qz������\ ܁�g��x[<�פ�?V��
��<��Z���Ssm�0����9Y�' )1��4������s��adp_nz��C�gp�$�����8�4!��C�M-����]�d
��}�xI�>����iU���s�p�����')���V6���Fs`�@��m��v�
�dߝFjO,8��}M����EW����f���/��
�t��nRC2��T�ʁZ�W �S�V"�$#
�q�3�(#��n�Z'�S��:%N��thϣNd�>\�ZEC�V����<��u��V<e$'�5
4�?�0�4`��bmB-���]�lQ:MՎ���G
��ש꺥Vנާ�I{!Ya_�L���*��b��,�B:�VI	09���5���Q���1�4%�lr	0NjM+Nbj��?�!h/Ĥ�9[�����ʙ�2�O�Z�z�\ ����� �6P֧u�����O��wO̖Pڵ��^m(�7�5�4/���A}-&֚�ɉ}t���r.��Qf�\���W���<���,x����)��{�2�oW��t��5B�ඃ��C�g�5�T�У?��`�gx��s��\�N�sj%ZL�j��]���hJ��F����'����H!�	4����t����w$M"�W�+d"i�L���ok��������E�!bW]r��
��?1D �m��m���z~Rn��@T���-�c����}�XcSN���B�φ���G����e�����޸=��n �{�!�WT6�d���J���QM�B�~YW-4�0�O�]��)Z�3���N+�*7�h�"nz*���'�V7U�g������iݱjlu]�ݧԸ����W��3XE���	�:I��˷@�Z���x���u&��+G�oE�^P�!���b1�����qx�P�)�]�;w��_c!��<g���Y~f�iBپ���}�TS�������=)��m̆!�8,�.!�VD�P��K_��!OX��2?Ce�҄������M�����v�.%���e�a�6����䟓D��8�i�%T"V5u���+�E0Ko4�v��
e)�r��r���v�h���'Ѩ��$$��������7��aT>�źj^�����O��{3��xK�4��$|��yc�<���3��U�w�6�2/�]K1C2�2Im���Qu�[qx}'�����?<�cw%\��&�ضm�Y�m۶+X��Tl۶͊Y����>g������1��g�mN��'QIkOU����4�g�l�W��E�1��*���|�����;ܯ�7_�U��-|+�K%jU��f�H2����i��U,q�ƨ�nO�U�I{��j�BBwU5?�Ѡ��tB��ɉg�Jr�{���wL�.3�-GE.j�?��ך �Vű����N���M��I#��}&�<���(U~�4����)���:�;���Mߞ��K[x6�jh_c�5
'
��
ߡr�jW`U6�fLm�g�n��6e�����Qp�mm��iJ|�	|�'~���>�	����¸ݦs|HD���n���!��yG,y���*Gu��C��7�y@f@c�B��x�XU9��Y������Wuަ�T̉���D�}MD��*�?75qT�WBE���ld�c�|��I��n��澂5wxCH�:d���u�SyE*bPI6�9�{Ϊ����x�W�ݭ3cݥl�`DR��2RQ��k�w�V�Dw��n�v�n>]���Ҽ|�h+��PCQ ���.����[4�/h����'4etaIbl��1&�'��RH�0d���'*�^:�{gN��>�\/n��+�T�`�!|�	��"��lTd<�N˭����"��}��`�#����m�� e�r^���0�_ݜ!�`ԅ�b�W>�]�o�0��K4<���]��|��}�y]�Ј>Q|OK�_m=]Ƃ���42�H������\7}��Z���Q�T
j��񮷷(�*��4h���XL���8j Vբ��Pzӵ\χ�p��g>D��d���U<���>S��L\{{�Ŷmm���Lu��&h��<1-��A��Q޹�#�*�?p��ag9t��YbpR���ydf&��fGU��}�y���bC��qϐ���_�������\l>y[Ӣq�p#���^���p'h���0�A��~iqs���mk�/A~�4ߛ����'�\����d����x��s��҄��O��]�ZGi�N	���%��h)����-^�<����j���6ͷ(�p�O�R~H�.�/d-Y^*�Kp�4jEu�JW|>ߔ����a���H�<��A��zF���	���(���M����� ���ґ�?�*�/e����Y3}m����ʺ��$�Ьs��$����D�t�k�Q�/,�qT�M�l����������?�y��h���˗�U��B����bQj)���d9�z�G��˧xmd�A�ZM\�,�8�48 Eu4�ޘ��Q|b�'�+4j�'\��7W�c�n�o��RkDu*�n�����eY��^����c���3��,���b������.��"�vf�C�ZnMCR�U͇MjvNٳ��p���˛��<��I$�d;��&	dDZ�`�Q�"�SF�ߎ�
]���K�^����9�qQO����M2��«�_!;������ 9�'�I�(��G�rw�$4�V��jRy"y0�Ӌ�'ř�?��	�i;��>UBMO%�X�#	fh2"%y�'�և�T�9fk�ּ�!-O�)��['^���<~�h
�]��u�q��%�R2+��I*��%s{��r��&��y���Ӯ��8����"S|�GN��bKkӐ���r�BK�Y�a։Y�X[|Vh-ݭ�����I�BSxo&�5�]gS�Y/���b����BƆ�N����nG��/�����|��*G| ���=�7��x��(]�4¥�v�ɳj�Yp���d5������Uk�)W��׹���_�I�r��6i[�L��:V�>��H��R��*Wpd����a��\��Gv�д�Q��v�L"R������Д���2[\s��	�R�?<�<��"WK��h�k��{l������k�����-� ����Q(��	γ$9����̍×m˘�����X��0��e�R����u8U�,1���D-[ΒE�j`+7-Fe���U��I�NI�e���V�i2x��a�x�o۪ki5�G־�a��џ�o������V��h���8%��Dcdl����Sv��tn�zY���U������~̯���Yc���s�+���^�;��� y�#L��ꯨL(&i��YC�������u�~A7 �l"�(1��?��������x� ���e$��/iS�"�8�\��2̈��=�&/��K�s0Sc���4�a��%�b��`�m�Jy�̪��M�U+q��(�C�G���4����&o~�L��þ\�M�B����GWuMu�;�ri��� ��CGj8�o��J��}�ʱ{�~��v�=�:H"�c�L�v�XXw���~m�ͩ����	M*ZV.��K�Mx�5��F����C:���3"��Ue���h���ޅ�[_��E]�"ߴ�8\�� �ȭ+��~�_�X\LJH�5�sؤ�Q�z�q.�L}_�6_�v���K�r��Y�P+P�Sws��z�~��M|V�q���[�	�����	�V3*�84�I$]��xvL+F�ς5�L*.�͆8����qj���0���4Q�A�$��(�5C��̥F$W9t�<���GA�|Y|�`=��H�"��9ȗ۞|
���X�.I�$� �+�\8��9F���b=*RbeU6Wn�Em��%R����gA��hϕ�_��h�7����b��8q����tX���vt<gU*Ԑi��~j���p&3�G��h�2I�� /&w���%����G1��멥� 	��S���^��o������bl��QB�E�<�!�0�~�.NF ��A}\.X[�4�id�x��w07)�Hu�PHRu:��;����	-��+��=�3��\�&~��� �D�j����d��5zT{�Q��(%�Lv{V.���-��DI���1"Soo�g\���O�[O[Ӷ�j~^IJ���������'2`^o��Az����a��^w�%Y�ۨ.}�'��q�2t�zM�Z�w�����
f�՜�(#ñ���[5 �6��f��?F����/u�غ���V�C�G��"�ɩȤ�zC�����7:��I���R���)��st]���B.�T!i��^tg�J��V�U'5I���_>C<�n���Ō���Y|��`�"��^�'.6�/�u�VⒾ6-c�����m���W�G�X�����G!zeE=�\�m�9�8��M�${/G���-��Q�
zO*ʨH�8HϽ�ˬ��xdƠ�T�j�5�ѷ���U* �G�*��`���֮]�b/W+�:��S;)o>������bLl��,�*�l���
��F��,	fḛ����%%�OiٺC�KU��P���r�� wf���bŰ� � ��HS2t� .�2�ڿ�����ky�1}���k�B2\@�[s�)�y�����}@Nyg"��u�	]����F���:�V�������[4�gR!G��zT���5����Sj�Y֗�s]H�ۛzʏczGݢG]��c��VL��gԚV��'����הU�Ă�i�[�:�);u��Z��p�Z%�
�]�3��%iľ?ꏄ��c�Rj�y+�8�I$�J�u�d����~=�8���-��>��Ҷwgi�T�n	��=ii�/ƌ�/M3ڕq�5y=���]v|8�><.�]�{�x�|��3�L{Ȩ6���V* l���_��{.��BB�㠃�P�gͲ�oYZh�+6�(Փ93�Q.���̙U�I�B���nav?�8k�e(4�!=��/F!=$e��<<g�$�+�;�u�iǨ��o�G���K�"s����WK��� ]���
)����7p%pg8��g��~߱n.� '�y+�^D��:�a�h�lɄ�}�����ƃ;չP�Vc�]f9?+R��	9���h�0���O7<
�N=*��aÀxS�!K=�Ai�3�YH`?���U��$�g�30���lA�4����`]	�;4�39�Sh��oI���`��������6�"��_��d��oiZ<��)���U����mm*'c1����\�4Zj���jz�wz��ysrv�=�Z#u�զ1�Ն	'�b{��;����菚?P-��R%/zc���:�Gzg^}�Nl���˦2�yz��x
�+����w]ߖ�_d{��l��ŝE��-����&Bz<JO�(8#o�-��<����N#�}sܯG#�r���&�ͦ�F�r�:���w�B�A5��_G�R9��y�e�qw��mu�� ���+8��L��q=��{�c�?�0:<��`:R�=����Zr�(�Jٻ]b�4%�4�����;o���>�KJ������Oy�Arp_�#
�r�p;6���.>y4I�B80/�3ga�xxG_y�{����ڴlQL����*�E�)�	 �B�(�v|?�ۢ�`{�D�xE��pD	����U�B��O�N`�v�4d:�N �L���|1_"����M�ß�dA�CnC�^T�v�{Z����Q�C��+���Ts7Lf�}��������9��a���1��eX@D,�\AebB4���uϧE�"H�{
G)�)H ��p6��#L,�nTK��}3Q~�-��.�H�/�RG��k���4w߮���>�V_��MС���k�����֋��/�С�x/yT����<���#��"��l�Y�׽�����V�T�q�9��7��$Z��u5������&c�*&G��fg��E �)���j�S�1�Η`9�d�%o����N�w� ��r�]�sG�����e.�˙X�-�)��\a` �;_�x:��!5X�8�~$X��Ȟ�	WȨ0�C��t,�6�a��Z�;@��6�2������m�.�|�	Mi��W�=�:N�6��L���T�b����{��@j�!�����U�Pm[-�D>4���D}j�p9��ī��s`)f�74����L|��hn��)Nв��~�L@�=�'��qߵ,l}�4Q�wNg�js�j���k��z`sɏm��%.���Hp�hpg�IƷ4�����ՆX�w��>3���њ#�şTM_�pM���fNX=71����d�ɋ��W��w��h6ͷ^c��X���F�լ��Bs��<����v�k��<����m*P��TM/�jɁ�@b]ۆ��bۣ��C,E����M� <���e|�֏�U�4$�Ӝ��a�j�hT��e��/��& �)3���϶bb��	�,\��=im�ޣ�dM�8W%��gWu�3yǙ� ۢ��_���}g���u�M)߄2-Kn��\��W�m��n����8k�X9��J9�!���|@;���~z��nc�$�O���K��U�ۡ�o^�kv�_+�k&R�3됫gd���1ehޘӦ`:�;� �����~J(����s��0�`�&I�1jЂ��?�5	��MK�.�c$d�Scnm`�[�<C8yH$P%�%r���r��g�zg�i7�R���4�����j)���0cA�������jk��CU"&	��i�]��0?)��K����|��]��F�~�^�h]����(z��dn���Εz�O�@�۳Ha�����%v�v�[�����'�YDY���[SH
�E� yK$cIj~㆑Z.�/�8�Y�G�v%Yl�2]���zV�FK�$c]�H��G>�/U���"k���	�m�G4�Xu6�#-T���LM�)/'�ǵ��1J�W]|�KW�=9��2I�.V�?<�P��<����qj�`���0qi>Ƅn��2��
�@��TB�G��aE�/��9"%{DX����Z�u�6q'iućy�E�h.%�w�Ȟ��B��{��F/�u.�݅~�^��L������0�#+9hE`�(���ʲN6qO,��5x��O�~vn�B�>%�K�;��ް���ovD�jwl��RȏF�L#��r���ݏi�f�����4�#K�G�⫔��U�?و�KV茺�N��-i����!V�p��԰�cb�qV��W,Ö��o��R]T�z���kwgh��Eh���r	!c�e�%�Jڷ�b�v�ς�"���������ŰG�"@G���8̐��\]d��V�y���|/��h���E����'C�k)�X]j&�(�cw� ���*>y�&w���E͐.�r��.ꁀ5+��U!���P�*�����>7Ĩ��3��5��������mL�]��������K�n5���݅ow�4xε3<V�4�U���=A�f����6��5��ՀՌ!�c{��"���\tX��^%��I�b�ѸiL�x�^��f�8�񋞝�MX!�o�X`	L����.:��9�J����߄�ih�7&��oA������KH�����jT�*�	�P�+�LK,�� �H��̔�G��Ad<���	�z� ��_�@���5��+�v:��_��8*���i6mk�Z#�\Q����'<��4�1đ�[M!��;�b�|�w\�kG�&=#�����lb�nyd�Z��܃608��5m܏���Gs�)pSSr�Fy��S�6lV$�����-k}�24`�K������|Ř��&ʈ&�>Zv�R��b�L)��b��x#����BLS��3�7�R�'��,4��q�@")�� (���'(����o�5ҋ��0�
D�rԤ�ï�[�?�q�%��$�x��&�s����@$�Ÿ]��I/h#ٲ/b\v��E𗐰*8)àsc�C�`ү�Ƌ8t"�:��̲���f� ;�-�k���QB�0�lAN�8���Y!���0����æ-N��m��#�t�2�He���f��8v�k�.q�/�PA�"��' ��_��8o5���n�8Cڈ]f�`� �Հ�m,k��l	؃�o	��c���ݔ��arJШ��J��p�����'��� ڼ>�Wle�a$T]��$�j��1ǩ����Xi"�Õ�U>;Ɗ{ n��^e~Nq�<K��+T�"�{8S9.��I��S3��͚`��m��ZhT�4ՠ-־Z��d\}��~�������vj����W��S]c��S�:�F�cj͙5?��� F��Ӹ����|�p7a�s��L��uG��W�Pu[�#�z7<nW��*�"A�Jh�]W�Z\ނ玦�Θ�!�nhkt�wz�Y
�]p�$��ʎ3HYB�:���9�þ�gc)�f�C��@�7���S�r��.�D�nB�2�'`���ߙ\��ZB}�	�-`��S^��㌌�2��Ţ�"�|ve�!⠰&��|��sw�f�Y֫E��
rQ�m~�Пq_0v����-U�6E����*��*kz�	ɡ���6�	�*��]��l�K^�"F��VB#ϲ�GFӖPKT�޶Ъ��ٱ2r��Q�_���E'^Q���/�B]�<�Ԭ���s4f�=���!n4�n|x�	Z�&S�W^�eA���]ŵdV��B%�&�u��?��0�������Y����.6�ݘ[{��0��tC�RU׿¶�c�5��a�����WH\�n���1}�V	A��mG|���M�WF�t��hHoDV�7�5'k,�C����Es��L��(�1�w��FM�2�ahI`��^�us\�9X�?ϊ�_e>�̡�l"�����~K��S�*��-��!wX8tN��s�4K��N[��zE�	�#���&&J��<lq֖R��Y��Ȅ��`J��D=Ȧ������t7�Zz�;s�NǬ�u(�+�,5��,��Eף���
�z��8}Q�����+�-�2�3��W�N��FR��\6�u%ck{ sL��q?M�ρ)��X4�$�-��\��������	�Vʡ[Ȧ�=����i�}��{ï�E��4�ҖM�ODܚ!�D��!X"x��_��;PȬ|-�I:��1��,J�i:�3��1Z�#�-�a,z!�~c�g�������@L��>}��A�o=�]����`�
rV%���ǫ�����Տ��먗��:��;�u�H	b
H��h����h���v��f��I��U3�B.���R��3�(�f�RX�sSeh�.�dzx�>��/!��qUX>.H��5�H$q�nx1s��놫�"�.�F�k�b��f��kzd�F$�Sc%E��:�'��K�uJ,@��3��ѼW��DX�ĳ�?{_d����f��Ĳ:7��.BҤ���p�0n7ɇ1MJI�`Ih.��6F�'�JbǺ !�Me,�f�"���,�+hF`�|����?Z�uf��覧�IC���'��͝�NI2�ƩÑ��������$1̤Fc`���̛��`W~*��[�xP��oR�b������b ���b�������!����%��s�(zۻq.�Ͼ�v�l:�����:�I�1Ƴ�b����a���ޡk~��b6�l.�DE��:���B��D�jQCK{
T��g�
��fл �QŤ|��re$��l�׻�ҕv�I'�d���Nv*4�x˞�C`h��g�菜M�u����o���n�3l�TzF��\��֭�*w%�%���c�TTFFp�Yt��h����<MQ�i=�g }8Z��?�5)ӆ�p�j�S� 7)��U\#��\��m��
p��xty�2���kG��E:Ju�!�U���H	"�tk�I�֐� d`�.�GQ�OkvZ������&D+����p�@�Iꠤ,�'�GRJ�)�F���+�\JdT�_�v��:����>qr$
����mk,����NA$���6m��-�|>0�x�m��%��>q�z��,pVt"��[;�[��LՅxrW��W[ޏ��W�[�C�Y���SH�Cd(J׬�Z��W;|o6�͟?�?�|�<w�F�٨���9ԋT�HSH�X�Y~�D�ߪ\��a���D<�$C�)+$�D�}�Aa��(8���O�{�1��a��p�r�&���Ftd��`@cW��ᅸ��uS*�VH�)\�\횳���h�kA�U"�
�����C��7m��V�����Z���6Ln�}� �* k��i���'�&d�/��O�5���%���G���$����	I}2�	�1^sG�Ӊܗ0D~�ڿ�|���P��C>�&8���n#��_��Qy.�h2-��tè�g̥�i9�`�=�x�W��<yi���v�Sp�mjn`�����G��3�� 	�]����_���ć5o��$���*I����*m�A�A���;��V���RدP�r2eb�USZ�s�kԶ�?.�;��v}b66�Y�x޿��_流�'�P]�^�w�����tƯa�Ҭ70Uh'�O��B�qRQD"ʤ�ӎE���������?�x
NW�ٞ��*��-㨸N��}Թ��ٴ���\�@Z�[jE�«��j魻
|�їw4O�����dM
Z&�OE����I�������Dyq��:�ی@J�&P]�{ጛ��H9��|p�%��]�ۉP�gIt>&_:e�W�7-E�P	 �D>{뙑YHhj�"IE�B�"�4T)��3/^�w�묹�:�'��\P�&>	b�J�w��������e>h��������ƴ�j.騻��v��Yt)�⦺ګ�J�95�S�-�Exd�P�4�v�Y���^���y�w|�/).Z��a��!覦��j���-@D��Mv������#r]����*����FUq�B��:L�[�>`�B�Do��A�	z1a5r��Yxl�{�0#	8	!	<"2��v~�����&d":r�=r+�Wh�M��r2�`K��=����A�p��C� 5���n2��-���Vh/lm�Hs�071���
(T������f �fЃV9֧
�|��u��4�`��V��%�
���b*�$f���̵^�B��L�Y��IJ�j��,�~�4�Z�!��#Q�9�����u§��/����IX�]��SM1G��n�����C�AAѮ����P��y�m,NҲ��\���βD�>RC$K�P)�9p�%0fE=G�l¢�b�W��XZ�������ǂ���S!�)�8�̖�t4.�|��2������O��_E�R�����T�QGY^��Oݤ|�O�W�ɥ��I�l�Ɔ��I30��s�A $3�0���s7%��Bt�4̆��|��;�y{�P7�Bߞ�%�J����}�?�hT
	'8t���7�IHHD  (���pЗo�q���N�M����4�߼�2�+�1_��@�N�����e*ٱ�=4�%�^F���=�"�C`��&ȭZ�W���ɕ��:�Tw�[�����fw���z��_��Eѯ\E�x�I�Ī����w��g�g�)����<*-)�/�kˋ�y^�o�p��ԉ (;	��V_��W�RYѦ�,\@i����8iݼ$U��^�v
��}q���l�u�s�F�(��Nw���I����((L`�X����:l^�*�z�+��0�Eo�)V�6�WVF�V!�c�;H�2p{�a8]�~#z1�~H	1P:g��]fg�����i:��:�w`�=^�I��aKj��X��+S0�w�����J�	���ܯ�:��v�{��q�^�4KW��P���!�Ɍ3��و)�
s�0�~�V�L՗`�3@�mhu
���S	���{E��_�~�͌�����
�8�R)�74ͺ� S�[�5r�8Hغ'#��G�xc�ٲeL���sou�O�?B�7fk�y�߽h�<�/W1����DH�����]��J̤K��9t�tfV��k6GU��g���<��� d�
�(M(��I"b��~�����<ǻ�S��4�U.���k�����������_�v�Xd���f�1�Rm�1�6�l�/��L��,�,����Wzd*�HqM���̂J9ȃ�A�L�wuL�'Ē���t�mZ�����Q�_��Q������+����L��k���0�aA�0`��/,��t��JU4)�=i�*U*��F��(��/��Е\g o</�L�n�-�-��m����ܻ�2�^!.�Td�)� �>�8"V��D���7Ԣ�E��}��H�i����[����+�>�S�}J>���W�=�%��s�'�\����5��T����gJ��\�]�������M�a�ini���x���L�n�zҙ��4��+���3������6���C���NH��i!<�����5����P��XSZS}�J����gx�\����3���z��)U�-*ǘ'8� ���0��:W#
�TWRW�l�7$�D��\�<�>/��u��	zj�i�^ �V�[+��vD�~�*��e,--�R�>A�:1!�'�כ��tp�3%�}�6�!�u�kg�nL�(��U6s�%E�������Ȅ�Rd��n�0co�?��.��^yD?�0
�����FJ�ŇF%Y��@��oC�2R������E�Wވ:����ⱥ��e;����u��*�f�6�����+���e,�6�c�.ѫ@�JQ���5'ȑ���o:@���"�L~wp9D��tHV��[�z���S(H�G$���.z���dQt�V�0�S��#i�[�]Q��*�'J����6����_kG[�������z��?������h��V���I�W�].�N[��}>>�4{gS�!�kJ�~ɑSx᪮1#�-k��s�s\��V�,�/�$~�P&-��y�[��de�ZRe3��F���#4w��D���}��D�8\�H���Ɲ\��1OV�(����=����ϓ��=��������w1%���C���a�M+��=6����7�W�6�c��P� �EXP?2>��1k��f'/���-��xc����*�y�p��l��-���N�CC$��U�Y}��/��4*p�/m'��`Ri��E~��h�F}�:�	l�. �p�Җ|Bt�V��T�¢kگ�x�'������)���A.���6U�l([g���Fblj�t>���>�:�yۮ��EJnj���D�	�Z�3����xj"4i�E����?��^�~�w��~+��/'+&��̃w�Y�G]�5��X+��O}��Og6��vȱ��^�����EtZ�}��[B�}�-��������v����a�h���~=��蕺f^�^̏�[T�̫���0���L�7��޹u�9@Ed�{[	�����%t��,��tT�Q*Mk�(-A�8�����T����O����������~3�����wo�}'kx<��boue�&P�4-����!�E�Qbx�/�[w"�o5�1��?K��|���pA�m�$5R��������y%8Ƞ�5������a;��}�2�;���Y�%XҴ��-�b���8��
�.��[�x���n}��	��{;��W���Tj��2� �+�t�'0.�|�U��
�U��ѭ���h!/���f�8�rʅ���C�1 �ք^c_�AP�dâ"����=TD���G�M���SFq*�����Y��M��diľW�lN��pB��������W����&�Cf� �`r�\��Lhch��r�ȭ}��h��Q����r&����ƋruF�p+r)�B���֮�*�on<(>�샃�����h�n�D3�(�3�JD�����ܵ3�,�$2�:e��v���<��}x�L����?9�#�%U��in��E9贯�j�����e��*:C��Sӟ�b�<z7m�0�s)��/����N3zxG���=Z$ZtJ2�����񀅉p�3��ѩge�X)����'���N�)0��j��>��Z�K��'�L����lML<@�����6��x\S��+*@$dcC�R&ojȒ8L����,S:Z�W��6�\ǩsC�V�S���&Jl4�Ԛ�i����b^_S$6B���1;��U-L5���Z_�T�+��Z�z(B����wV*ƽWA;r�/?��Kv�������ޠS�I�?3i�Gy����">8�g�lH�
%�������X�YY�I��ע���2I�Eϻ�T���Qg����M<�GB��hj�xO�;/�>�W���QZX����9�j����l�����R��ߏ�0����ra���d�����a?\����E�o+|���?){]]�kѡ�7��/�D6�t8JT�A�LC��\�&�6��$�B�+��߭�2CZ����(��d�K��yRea~1(�b�� ����S�Fj�kw�;��>���zwY���&n�{L�jJnb̫��w���W s������N�1� ݐ NB�#=��;��DEs|���KD��׵�j��M��?u(7�`D�F]�\�<17�2���t1Ϭȩ3���zЊ���*fZ������r�ߩJf��>� �&R����&�����d���p�o.�4|>�c���?�Eh.O_%c��ANA��#*�a��M�����A���[�c�;�S�Mh���)�^���<���кvV���6O�Z|�]$�y Ahi��B<\���1�@��<Ow�*�~�g=����c�{���놜�U�g�v���m���%x��߆\l���Uh�	�Xif�XhGϿT�%4u���ǽ�m�����[˟����D�C��}?aKd�V���#��� $�bf8�7=��G���߾HOOs�����R]�%���O`K��M}���W���zBb/x߮��f�ΠU����B�W�yyP�G��(���q�Р����c}J"l��������#W��#�;Ƃo/KK�B�U�<9qׂQ��e���jRp�*��
��ga��l�p��N�����؊P�nr	���ҽ��Yx��h�dSdՋ�ع���K���A�$�O���T�ѥ8G@�7&�+Kh��㯯	C�59$ue�ï7%��o�_(1e��Q`GkA��Vh��lm6I��9v�~���eI�P%[S����J2[C����b�z呍�1�g�p����N@la�ȓP<.���j��Y��U+�Y�I�V����Ŋ���nu�-�\���`�3�>5|}��>����~�q늖PP�Ϣ�T�9�4��ڪVF��l!�FL ��\eJP��EPs�7Q}�UP��G��  �ڒ#O��}�@��i�H	�ԓ��Ȱ�J�n�D����鸅$h׽Yݷ=��hJ��\�Y���<���-��N{6ܐ����@dD��x-��7M/ H�2��������c�x=7Tnʉ'����z����#�Gl��~���qغX�U� ���jb־���m�r����n�X� P�:dV�;#dU\���s�;���!s�����G,�iq���g�JkJb����,\��m�g���T�dv\�%'�yF�6g�r�`���3��bD�?5%�����z[���{�:����i1�a@���V�T�gc#��r*y�A��Y���L�L��)�6��#i��T��Ј�^~m�:bI"��*~g��)e��3���MSE�������%6����%ʈQo	�U]��Qxg��盽�2�. =l}��2M�~�`Q���EjΒ�����5<��K��g�;�|l�����#��ȳ��?�ۯ4��������F��������
���Ҟmh0�r��3�J)R�I�`I��QjU�*�%~qD~7[zx�l�����-~�D�U�9k�1�G�).Q	�����H��
*G:,:�R���Lw?T���l�F�&y�'��8�&v���nv?9���ژ� ��xj2zsd�(p�j�rKb<zC��z���`��� ����:w���띧y(�Ӡ-�p��)��D�_j��؝]J�M��-v�oh�J��'�N���YǚG>"0���k]��L��a�����5B˩R�#���4Z�"��N����-k���E	j��sL��y���s��\��c�t�@체��s4�^��Z���Aӛ���o(��i�x�7��O�}%p��<4��������c,�*�7r	�kkt����< [N!�h���Р�aӶ��F�\��������EVZ�D�D�� ����<�ޜ�T_��db�W^��޿և&�4s������N�0*�a�s�Aa��V�z�F#�5S�$�.W}һ����4��?276bM�3!ǈU*Ju|R4i:�G�yV�Lot��ߐv��K�o�_3���^@�u1MN^�V��i��on������W:(��q���DI������}�P��A�$l�pn�[����ЃH��vS��;����S�6�&�5���8V���3���^s!/���?W����&8�n���ȝ���R)���wt���I�k%y3"5��0�,��������Sq3��OLwM��&~�����w��	��5[�M�D�
�T�v]U!PD~���%�S>�^y�+��S3�Lfڻ�b��xL���*A����g��Xzc$��w�D�A0����`)S��.d)�t�Ht�Q&�WOQ���
��8y�v��X}N�������.G�W|�WǟT�y�d�Q�~u�;�Q<�6��}�<ԣ�8| ��	p�,m$:��5U4&>~1M��{{N���wP5��� TC����T�K��6�o肔8x�y�E�c4-�`�Ҟ�RS�^�K�{D�m
-F������d9�3�)�� �0�����P�x��1Y`�k��_�z��Y�]_�fs� a��M����;��tOSe"�n��:��_;�W�&|��������+���(��@͍z�V~<���ޘ]�N�V��a��5��c�B��!�J����������@)0�����D(x��>G^�R��P�0�<m��[�x
!G�1i���/s����J����u� t�W4�ޖ���������ܖy��I��~n�Ak��D�f�����s�g*��9f��Q'�F��d��C忣wy^��ܚ~M�g���KB�*�HH��A�DR�~]��/q�{�m��5����:��%�!b���\*>�[�nȯ�z�������/����_��>�":1%�"�Tȳ�
ȳ)#&��2;I����� � �.�$U�2=St�k۵���"�L�6g��e�@�7i�~�VS�	>\.2bfƚ�w���oW�A���K�!�t�B�t 9H��y��L	X�K��q�0rM��E�}d�E'G:]t^���|;��꼮�O�fR��ք@)���7���;���P�*T� Z�=� �k]u��P��-�k{��I�vf1��b�\=d�ϙ ��6�rY!�QD5)��g����E@N���7���^yLz���W�����l����ҁ�I5i�
�Fk�2#O]�&�&\cc���'���4���+	üwYU�d�w#П��O�|�J���O���́U �I��ƿ�^x�&��^,Xly�6��5�������(`�1?��s��{��))����r�Y5��>��Q��Qm>a�oK)���VJ!Hq� E�Kq	�ZJ�R�!�$4�+�^4��wד�9�y��~H>DV�\3����=w�I�z5b4t�T��1D��g9W@��������W�I�Y�[�^ۤ��ͮ�x&����j'c�f<����f�C��礡f� Q�&Ͱo�r��0
�è�=���
g�w	^an��*Lh�:�踓>��L�˃�D��h�1�#�z������೺1�nW*���j��7���?,�UA
�0(��M�Z@Vg��֝�5�z0:�m���p��������9ܟ<3cc0�7C�͙\�}�O�4��H,􇏵{4,�����6O��_:���?͵�>^�w����AHoY�Q���6��p��G�*�����b/W�W�����`uV5o�o�Γ�GG�6�+�kQ�OY+���"=��b�q���W�b�ܗ�^"�O��[�Oԟ�e9;'�b=l�4�e���od$�i���V�7�1��Bu��9B_�}����¸m���} ��AZ�mi�U����*�}>��4���_��M���#�"�l�`K��N� 'ƺ����K�?�g�X�r�§������)N�y�4���Q]����uT�-��oU������g�����o/D�S�n�!��-��8 $N�8�g�X��4�n����Q��	�-R��X}�$fm��d���xڎ��'�<�X�ɡ��F�s6�u��Pi����>���W�AOt�OqO�ijq�3uV��ژ��O�7O�r���L�DP5������8��ӈ�K7?�]��P{�d�Jũ�h����_��p�CtH�J���}L�Ip�[<~��Rv��7��hyxyE�)�Zb�v8,9� [����Cͨv�"�vv������ú*�' ��d�z�8�����&ң��v<�Nn$���QY�u���� 5���	Y�c]1)�|�k7x81��4�}������qU�o���)ȥ��迨j������E���Z'`�k$����5�Ϟ_�Q��DTq�o�ڑ*�_i[�R���"�m���%�7O��'�d�0g��@D�n�:;��dQ��p�m��U]k�0�z#�����6�^�%���u��k�wpx����W(�4�`X{�!v���H���}�x;���tuR�K���Iq�a��#weV�=i�g�ot*D���.]����6�r(�Z��eed��,��_g�I��<���X8ǫ���G�b*.V�Y���:��]~(C���G�DX�)��ǳ�d;&BJ���x�+�����__�L�N�t� ���w�ֺ��-���̢��Fe���J�O�>a��\����}P�d������!�}ik�A�,0�D���	�7gT�>�Qhq1�L�������l���M���A�S�.u��c����|�T�^�����dG�1>b�WBB$��xgR�0Z�Ng�.Vg�/�?���7�a�K�~��i �_
���`��%)�&�e���a�iڜ�Ћ��24��,)6|�0́$�;�`|z��˃��Ҙ�C��Ԣ]��;�U�>�s��l�ĚK��=Uѻ1��L:@���PVW��h�����8��,����bF 7��r�XB��-��FFq��>l��3f+�	�]k�sژJ�EPLL�Wzz{3rrz\��ED(����'��M;�(�q^ֻ?e�_�v9\��0������۷���w�:�* Cb��l�8|>�්+�a��?�Mm+O|娶HG4��i�{1)���R�ar��1p��i��񷶶��Q�Xlo��j)���	YN����8 >>�64�4O>::��\���X��߷=�=�2��X��s^�'�~�֠1��q�^�YIR�`�$��q���\�Q���Hc�����s?:@��hu��L���(���;ʌ��X�K"���(�O�d��� t�#�U(Vlvc��(ޥ +�߷I�`dL� 5�g�͟Yo�� �����.9°b@[���Ey�7yK��.�E��8�����1�r�׭��	P�O#������Oo�rN$@�X,co	o�*�a���5�e����&�`�R�,�3X�S��j=�����'�۷[�U��I���N�Vor���EQ��B�3^���!_�����R�ysڼ	�1/ձHnX_�1�~�A`���7~1����n��~�B�_���B� ��4~F-�]8����e	$��ӿSʕE�g�g�a�7���ccL��,�,x?-F���;C�Ky}��u���#�Z�����n��gZ')�i�У�^�;)
��LPef��!�:����LTQn�S�#xO9���z�MJ��!&p菼��?�=�@H���k	/���~�w��<1{��I	��_E�pw'�2RI���� z[�ˏ������?��Dvvv�	����6ݒ�?sXvB��R�8��I��[96yg�s���,��3�S����3�-,,fbc��Eo�f��ί�WS�E>z�RvI���&1腧F�2p�_�f�ϒ��l/zj��Tg�mBJ��c(+m4��㜖��&?����B@���'��4r�6���m:����|�c����bC�����
ʠp�C:��|��XI�}i-��j�N��,���R#{x��k��n�
�y:5�(�ʒ�T�?�i�i�}5{��ٛ��k|q�-���� ۦM�ΨKz�Q+Jg�{r��K>G7�4�]^�MN��1����ŰI{��w�7�{���=:��'�>���3�u�����!��%Wb]뷹���O!{�֏"&��S��~�u�jAFHȭ��A��1ɩ�;6q�h�e$�v�&H��ӓR��$�I�{��Z㣘T�7�Q����):!��U1s�3x��H�qsC���"�xC�{1���;<,�-I*,˒?����ڥ8h�����m�=�^���A�R??Ƙ�Y\�&�o���^i��߼�`k��L�M����6T@Ŝ�H�*xdP���(����+�-@|�> U�EV���Q���G��{>9!���38��'w���p*�=�25,��5��dvC��T7sc�?����/ἒtM�<�����峨�s�g1Б{��{�!k��v�g�j�T�r����B� m�WK�;6W�e�Ԉ��C;����0BȡO����Q�jX���x&��]Q��me�b\�,�/�⳴��
�l�#��R-�X��q����P��wEl��dg����*�%���g��V)u���y�Ѕ˞�� ����\dR���w%��0�B�2����B�y��9 Յ���j 
��c�8���'���~�r7���UqXIp���m��TFj^_��l�����b���S��������\jQ%n]9
�P�
��sp$i,7��mTi��˰�"��0M��+Ž����
ƈ:7���L̝}��dhc#e��[JJs���]m+`Ml/�e��� �߿���;�~�m\�Ů�o9�8"ӹ�e��[J�B=�Sݠ�ܛ��'�F��A��s���
�*���^�ˠK�_��_�����qø���d>~./!����Z�As˫�E��o���z�h ə�+~�����b_�XX����Ra���CU��\;�E�@$7^��8�"��ӡJAA��#B��|U3<]�-�5uK��s�Q�bޡ�vk���t3�[�;�S4- ��ߟ9٢m�!��W(1k�z*-7��^�}�M��;>6J����1�:������477{xx��-]���Տ�"6��5+���e�fZ�CUQ�v���I@ �P=^Ȩ볒㟑�v:ԛ�Ŗ���Oo������h��#�I�Ku���#)d�A\X�=��/ �Vh�n��4��!���OI���:f:(-ݟ�|@N�Ly]��	�`LP܀A1��4,$8�E���@#ss�*�̑>�
qUOKz�}��&�@�4�`nYJ�|�\;���t�_�l��I7�p����&{
!���$Ŏ�σ��r�;�H��!U�#�U��{ �� ����XXTZ����:�7i�,��%V�)�9HE_�D�:��H�Fۆ�E�5�4ٴ�B_�J{�s���y�揽 8�7j����WI��S�����cw���6���\X��<#�,]M~�Wd��D�T`�H����'"��h��Ƙ�ͱ�/v��� R/�P�dca���D�^6�ϒ7���Ʃ"������t���ߔW���w5�������z�����W4+Z�A�\��}�-��o�,����d��T�P�Ѱ�:۱��� [�W�g�r��{�J�#<atD�.����$K��Q�׮�]���>>�[�9Nɧ#���J�L3�v��Nd�Lh۴D0���aZ%�ۛil�U�pC�^Q�P���!z���z�]�"��Km�	�*Y���� �C��^T�	y������p[�`*W�G��;r��)A�����Qy�I�)W\�P9�ڰ�u n�N�\��� H��z�_���N���'V�Z�Z��H���.L|����[~�&��+N�g�f�t�E�B�����1�t�/�oVg}.p�<���BN�*Z|�1HS�X����U�v�*��*��l�c;L!�x��ڠk1�(�~^q5^�1t.4�v����Љ��9N�2��nd``p=\K�H����=�8�'-���L��F����cd�h4f���ɼ�S��M������g���粺�k]l�:g��D[{��FG��Κ���q�ԍND�uIQfa.�)������y|4K��O�ʥ��բ��T�����7�_ɔ��[��S��}x�5�hI�\雌���'>J����w<'���l×)�K&�!Ϻ�]k���23���QDUX�m�b�)�Ϟ�/�1u���������U���d��;C�>�>p$�¥���+��w�k�êȸ��{��M'~�v��>c@>�7%�z�ʖB��Dj���)�A<_�l�������p���&\��EN2��X��gj��M�X����rO]�Y?�������T� �W񝡀�WD�����m{�5he>�ھ��tz{�<,�a6m�fu�w���m�l�X�72���q��	^�]:Wv�C"}���Ӿh�Ρ��u@*���1����-�8�
�:AQ޶��<�]n5b#���!����M���ۜbk�T�?����v�axs��h2:7տN�^�SM�A�RF����S�/��,a��%~c�m���w�V�����X��x_wZ{7�
z8�P�S�"��������_�g����35�^cMT��O���@U~�e�j�ї�QD��=��4�%/��q������h�d�sY�bƦ�>��%��%��v��+qҴ��>�l�6�h�w���rM �n�����wrb�̶p��A�k2����v���M���ot��ʀ"��W���*o�GF��[[H��q�RS5�"����Q�,�F���Q�
=��{�m� "�if;2��9�L�.{ʎ#�	_~�f
�#lnF�hl��0Ԁ��x�z���'�#=/d��� ��"��%��&9��JN�0��oJ�a08#L��������i#D��3}Tm�6�>Ss�� 6�J����YEm��ˊO�ZR�����tT�z�&�=����^��Ԕ5
g�WSçp��(�M����"<3�ӿ�<�y/�����S����g�?��M��*�[2�W��r��%c�r�hT�
��&�S�S����r%A�xsNp|��f��i</�7����<@*���sP\K��������l����.;Ш��<�F��r{"Ű�ǛV=B�}r}�;���r��v�v�uN^^^inA5�T�Ua�Q�tx���[����Vƥ�*�Z-��3�.�� QF��$V�=�sr7&��S���s4�������3�7���V��ϗY.��s�|L��t.qcMy���|���1�ѻ"ޚ��Y�$w���erojif��g�ɉ^�����RKQb1���ǣ�E�!rh��>'#㛏>�V��B�]����EA�sv��4Z�#�><3����8����|I݁<�Le9OT2w���
,y����Gڑ@W�UXRrx��`��O6z8vؿQ�q�4ܫȰ�g�%ƭ��TQ�/�Dae�5g �=߇=�a�kjb��R�C_׭L��򇞛���:��p���R���s�^ (ֶ9�s�,��p���֪�n�gf2�SQ�V�}|{�`�o�,\rqᙟ�W��|G�52;��r*W��Q�I���S�fi)���A"��Gq_nVf��ϻn�����7�[j���^�pX�	�Ҷ1���q�o��T1�{;����-�wñ?��7����g���� qD��D����,J�j/�P�ۨA�ڤ������&�����)u�� �W���9���F��ϧ1�F�CQ2�f�2�F!D�٤_vu hgo�Ф��[��ݵ�ݳA¶NJZ�d��S�5���.T,��<�1�u��������g~����Q�ZT�S�Y���8	�0i^q'Ȭ��RJ�c�JҲ�*�)<����t}���>;0���������$��
��6O�����\����H�1�_)_�
��#��'�.�(lc4BSlb�t<�.�~�x��v��� ��a...˹����jka9�$zT��S������${��pD��&"�l�|rЍ�������
����,-�,=�]'uIY�s�~���A*��*���;Wm	ZN�N�ݑ��i���ʽ���q8琹�[�����c�?�	�|��X"S4B�q,���#%�7'"�1��M�{�:3����&�S!�)|B|������n	Eo?s�;r|k�������+#J��G�d�G�"��e�J�f�M�j��v�(@Z˹$̮�_������ ( Ԃk��v���T>�,����H�l;x��ud�Φ#N��)(~�ٙZT`y/���kG�fK��i�$+��LJ�Y7�)�+�y�8C}TG��EG�N���T~����x�t"�j�I�Fl%�;��y���2 Ŕ:7�6(����B��"�~|�6e��`�
�Go�l��w�V�L ��Ύ>C�q�?U	"�t͔�@�`���Æ"��V��gg�xx�	@X2�'S�l��h�Q�.4��H��۝��j���U'Aa��:eHT0qT����q��:M�8?�[�|)?:XHʏ�t64�B�L]sȭ�RU��_�ޏ���Y�tK�q|�*��l���Bu��1ƌ�%�꾊�֓�J�]9j���k�`N5�X�HǀZ���I{{_͋2$��M�k����}��1�ww�W�~��d��H�T@|�V��8�<\��/�Qxc�`?� �C�X�h]DO�bA�d��Փe�:졝�E�������@R�ϔ�7g)�;����n�׷7]A\�Bl�YE�"t������O����f��?-'�c�8d��/RZ�d��rTQP~�)C�m|�B�h�����D�֍�'y.� h�Ly�mv�)���".ɛE{:�c=�����S�N�4����:��0#����F�	(m���5�38t<g�r?�����4��O��&���8�U� 
���vz�J�_>����"mC��@-���~�abH�^�Ī��-�<y�"F
{����+�kН�lL9��S��uh���e��2��"7)��t-uפ1i�OѴO׮ 㑱14��I)����0��Ad��ߦ��K�{�[�$g/��4��m��,�u<��K4�Ra��xx��(7[�E �s:@����;�,PVb ���PQ�hZzx�L���Y�k����������<�P��[�*-W�vZ�XS��%�����;N��:7	v'���]�ʦ�|�G�Ȩ�����p�BJњ�B��!�rS:r�O�!� A=�����|e�O��V��
$v.1H���q�s����7l�����gV��;fX����9�7�-tP�T���+����ݰ���`Gv��R4��L��W�+�7]͖[����N��G�����ΩV��d1f�����~����{�I^�̽�
UNA�������2FG��`��'G��y��Ǻ�b�����]������acP�t�e�����g���P)�Eiޜ�3#�I���y�4L�=É'��<=�\�����ȡ)u˖2Ho��q��e����
m�YS�{��1����on�m����I���f�hW����Ŝ�X�J���7Uֈ�6.H�ⷱ��!�����w�/�U�U�ueh(#8?n�2�r��q��̷%g[�$��#�4����a�	~���X���j�m��N��v���'��`T9�yT��y��$YI�b\���-�ɤ�Ӄ��,3,ϐ(+�����_Z���?��օ��w�\e�e��f 	=��H�cs��r�4;��~**Cm!�����&���=dS~�+a�2Q��k�-��%)T�	c�N��[[6��ݮ{�*�8�V�>K������O���'�����n�Ɩ�#f��~v3�|P�FR���=U,F�;�r�-XbDO�Uxw����:Bf���5�)�
�b�P�w�]��d �t�	�~ͱB��RFű6��Y��������wm�*c����v%�~*~��ˎ�ˢ�v'ظM��Mt}vÝ%EhY8J�W���z��Lý+R�E�e"A�4��\�l��������uZ���<2�Q.3h;�sOq͂q�G��ȅ���ɖ
T��-�Lfp�b���ۣq-0��@ۈ�âci��`��Q��#��1O1�hh��L9u�Ժ�*宅4�O`����$�������V=w��&	��w�M`���r�f��:,K�[��l����2��3^�%�$���l��ڑ7H�.>�99���E5%��Įm=b�m��:�]+�>�`��%+,���u�z�YZ�Us}�V�v�]��b�ڳ�YB���j@��k����ҁ9*��)Y�����W��\�`��e}G&*2yYu���=qg�|3��Z��������}�ТX��]�
���������yTiكw�S/Q$ɦ��ůip��d�&R0謶�-̌����G����d�����b���WdJ��:R2����a��1*ܰ�p�#F�)u$I?*�f�;��r���t�f����ܧ��pW��)rg��FC�քb\^9�����C�?�۷g�-/�����0())6*���<ƿ�Xb�����s�}1}�G;�Iv1b�N
'(���������f ���"���k���*�������������(gCg�<v�bC�B�`f�����$�#�j�V�0Na��uo�����U�ć}�{�I�^��0-y���X��Ҝֶ^\�{GȃEa���d��|uq�~��i��(����e���_{m�Fɴ�W��F��N��o������h�Q~)=��p��d��A������:�'����,E�� �����)9/��\{����Ǧ�	\��޶5������|��������%���3O@jS���D��(�'�O�'���q�$J�h޻�s�.C�b�ߙ�/j2ɱI1�������2�vz���Od���KcK�t<M�v6�	^h84����NMM��t�p�Wo�zq{{+-�=�1���jEӭ.�e�^6�bL��QS�s{{M�Dli�oR'Ӭ�{�7���ܑ��<�p��0\�=鵲�ɏ�Ɔ,<غ�x0� F�!89Ѻ*�H�<<�I�X�-���m�Y�Q��R��* �[��w� ��ե�Xx�:<�-$D�?"E���Y�J�y��1��ObG��������^I�A�h�ޚw�x�+5���	l���8��d�� ��O�͎�Ŵ�sFi�ǌD�BѥC׉��j^��%��Z��̣E=o���x�����=��T�σ8�5�ף骜d�g��Q�#i���^g�?WϘ�_�ċ��/Lc��t�
Ph��NN�;Q46p��H+����`J��D��ky��=�a�&%z�M���P5���3�����T��LMГxCC��@�vÔud�O�%�>����N�:��1�m��P�z�`�?k�Q�1���ۤ�����ߚ�����/��f�"d9�տ���8a ���Y�&�[~|�+��Ux�{�?2�\!�(MgEo+��r$�ʛ�DG����棬�V�w�����~h�/�E���䞁F݌r�o��6 "쓥�	�[ox.m�E"��+�T@'E��K�|j:�&�K��0���b��ϫ^v�Ș��ʧ'd�.ք���!ifK��Fƌ�_��?T��S��']?A�Lr
1h��bd;����CpH��yEo�-�����C��a���c��C�1�"E�5�)�1�R�$���{�$�Wx_(���I�lȷ�ll]~TT| �!yNp�>_MMK��^n46�a_MQC�-[q�ZC*̶䥆7�`�13�;.8��Gn��k��5��B(M���W�ΦR����ۯ�<�v�ކ�,422����(�����Z���7Ԅ��ş�ٲ�n��/����`������4Sp�A�#6Q�^��
�׆���P{�.���_*��K�82����⣇3w���߸�Z2n�C��J�!v���q����ͼW�2��Ғ���Rr�kIB��[�}�՝x�GI0��UN<��LTt�p�v�F�W��G��MȤ1�F#<b�O���W1P�b#�q����[e=�ތ����m�T���=�Y<8)��Ȼ��;
&"�E���&�M
��L���y4�.c"�m�b�p� �|�f�"�R�|���!Yz��J��d
(1��p��6��������J�J�E\�W�ir�ք_�?��x<��剕�_/�6�rf�2�HV�u�V�rو"���)F�뭳�CÃD��#e�T�c��E1<|����.F�2����k��t2y�p_��7b"<;sY�JJ86~�D��E���"E&7���kԶ�c�ܫ����ЊF��l�v/(��S�
���<=���W/�k��-�J@�g*�]�TF�� O���C
����q�SY'qԸ-?�WLy��E���@ю`�E�\�/=c�c�\��f�B���FK�)��~9qVr��37�^��3AC����~��X����+�|��g(��w�@��t�^ᩊ���z�Ҕ��V�1�T���.�Ej�RHD��e��7YM��v.��D��F��>L���9� �ttuO��&9H�b�@�_W��&�R��^�C��Ӯ�;;��+B��b�~B���(�N=c�������ҼJ.rj�����)��������o77�c;N�j�	/DEI�'sSS	��J�x��Z��&�"�"�ԓZXh��*���#��l�AI��0*����U(r̃Zgj:�!�}>�ه�]\\؈!p��j�2m���՛�M�O����U����Q,3��I'"�4��Y�B����.R�ͯ���,j�~���gZ|�;&�*����sjz�/� ��,gjJ� �*ӭ($�B��XP�\3	������������sGr�J@]�Tӳ��ܹ�]�>�h���=?[���HM[a�D��WMehfC	>zd)ѿ�
�҇w�&�?���	�U�~\Q*�Hiah��uf�re��I�X��mϐ��\����hQh6�A'*S����:on���o�����n�g"zG�Y����t����<F�A�ga#++�0Hʤ"��\{K�OxH�Y����}�2��uy+1�?�\��d�i��!~��c�G�����N*�e"��Sf�s�J��d�n�T��7�4;�W��iO���{���Ñ5U%C�|���/��s�kB��O��ܮ��n����n�
t��:GE����WW{��_ӹ ��7�I�^��s���cWpB�sj'Ԙ�a�o*�U�Ǘ���k�z�U:סM�`��>����Zr%��˙ �7��%�w
(�R��k���푅��O�l�hP�Ж� �O�Yx�p�(;����Aw2�(k@��t�`��&��Ym�������O	;� ���*1$�i����Y� Ldq����o)R0b�%��`;fo���F[Ά�L�j������u�����N���9�������O�Pڈ�׹m޿9����B���ƣ�R�أ�gΆ+���^b���z6bʾ��뭟�|��:E/������_�~#���+L{�u��qj�Ny�=q���Ќ����%�쾉Y����{�Ɨ��1^4���͉�#E�V��gU?���؜S��89�o_-\C��G;��'st�m�!u�6�>.t�$�J	d���(��w�����fX��"�W���/oC���S5BB��!�?�N��,��Z��H��@�U���{��H���}��s�V������_���+MJ�����@� ��U ��³ſ�	�6;���aw���qg�q.]����z��~�E�ٰ�����{�6;�O}��������������'����^U`��F؈�hҚ-ٍR���s�j�����<��۷�eeq��LDm69�����孹���l����e�uR��ٟ������G<�FYe:�R��K�+�ba�#�u,~4�Ǚ��6�X�а�s��G/`n:W*���?Xiæ./�/i7n�2�Z�>о�տw���CY������Δ�mwQ+=���`�+�B������o,a$c��x� a��o1�ye����o���E �&Q,M�T��V�A�x�j����y�����lx��������=��y^�핀�._i�[)�u���vZ	s��9�\-��Gk˄�5�a�=����� ��w;_f��%x�����ze�LJ@+
�o7��#�6�#�S&k�azVv�a9��^b�׼��]ՠ�}�N-)���g��)���K�ə>��>MhP-4���KYC���HYI}��@���+�-�\�z�My���W�~��Jՙ��ײ��z-�k�>u��C�r䩘�JĆF��ܟ4�ٳ�)�:�ͳ�ߠ�7�-��&�a��R�?}J����U�->6�Rg���q���|�Ȝ;��e�����g����^���*�_��t27Dl@Q�T�k"�=m���Z:�X<�C��7��:��̎.�u}�fD#�����O���u�LE�� @�C�a�!�6t��Ͱ�h^I��m�B>W}w/�_�b��ԍoa�h�U��,4\� R:����06��r	N���!k��܌!�ڦ�U��J�I�WXu5x8�I�2����ˏ�;����pV�J�֘G`�H|C�u�6W���$��B?�o�����5�D���ޑ
�Y>��������s�2�Hy!�G%���i[c�2�Y55>>��=?tp�x�1�fKq�scR�9޸�W���O]��?y��?�Pn�w��ƹ�uaC��:��˻X�\D��Bs	�ĉ�����Zwޫ�f���lF�gL0KA���?e�}H ���~���N�!���t�ڐ.U���r\�q��V���?��X�u� ��(O�u��{�z�����T���~l�����!�� ��/Ot�{��r~��	F��\W���a��כo��,WD�m��c�N���紱�<�U|��wVB|�d]��bד۸�<(>R��.�$%$�R�	��$��)���,�J
��1Z��8HF/J�?5�GA��X Ԍk92�`N���Qs�=�����o3ƝA�F2*ĺ���B�N�P�aD2�������ׯ4�Y��\MX"葷�����9[X���)��1�R�V+�L+�R"[6�L��%�	v�Z��#�;�T�<<m�q�����^SG�u�ͅ�Fu����/vN �`MR�� f�k9��>�||����t-q8��=�Ք�?(m,�9����"��B������m��ϾA��H	��=�pw�&)F}Wxld�8�C!�9m��Ƣ��aX�7�����x��B�n%?���]��''���x!�࿯�������M�ȢlK�ZtM}C�ޔ�75�7o�EZ1�k��n�+�R���.�D��?�j��.��WS�H�E�'�x���Ú��n�H:{�Ɖ{Q�y~��0�� ���sov�ra��|�����?宧������d�(���A^m�	y�;�X�ES�G�b!�4Z�zO��U��+O�X3=!n�p����3_��{lM���,����2�J���5�dkhow+&S�͆{�ՉO�Ӏ�6LcYs%�#]׻C�'��8��Nｯ{"������L�+�IE*�;Sv *.+ �7'?OUQfI��zXr��WV�����xҢ�;���`l��w>���>-��e�}s�������,��z9#t0�;��8���͆�r���4	�g��A���1a51_4z
0;20	���Q,}�	0_S��\�oʖ�N�{�/��<NI�B%��OY��a�����QFE汀[��n���6��;PָS��K���)H���(El��l]���1͠m�ḷ�@��Z��f�X""�;�!p�f�������G���l�X�А�J�o�I����>��i��a4J_�S���b�R3=�}�d�^��7��x��"3�Rc���`m�0͟|�Tc�$%,,,����[ן/k-����^��%��:4�ի���;�&{0�
O����>r���~���Y1���g�ݚ%_��������<W��ɾ�������?���W�4�_�#G����1p./$|^pu	lJ�d��9�8�����ȣ��i�~�W�7��#�j�?��%��`ت*������706~P�]<϶�FZ϶I`�:]���B<~�}z8k��1
"��l���I�,��xUd�vW�N����}�)#����O�h,/Ѱ1�Wi�7r�NI'�w׃6kk�e�6_]_��y#�'oΐq�w��T�B}�qbR����P����;��jt{w;��ڸ�X4l��^Zf�60�Ϳ�*�Xג�_�p���޿)�Ť$���m�&H�k���xϠ�b*���yb�]Pj}m���e����>)��5�㾞3��҄91$��R���2�I��3�/F8���*�;7:�V(q%?�o����t� �U�X� 3���JkF�?����|�Q�P�ma��f?�0	9l�~��O��0ɛ���D�c�L�S`�{�qK��l#���d28,�H���6tQ���74�V��gjBB����dnc��Im��F��IJٽ�����z�r�M9[-q�g�趙�̠�}L�zB	 yR�|��U��؀��֦Q
:�.|��a���|���K�d�\�?O$��E�*���-9�{��6�*���Ԍ�.�n^~�	����~c��"eN*��Y:=a*v6������ڃ��`K}#x����\�n�$W�O`�r�P{8�WU'�IL� 6[�8�J�:��b҄�~5���:?��*���k!��p�E�C� `Gٴ���UW�����n|�u;�Q�m��[��Ah&�a�'�2�k�݈�q��e]˷gK|v"�H�'�+N�X9�
�q��3�a�F�AÃ���<N��Dh�_>s�-��r!�O(�����0M��?�\�^�M�J"X�o��U��ni[X<���t�L�����0)V����1��7��J�Os=v��|�3�$����5c���:c91���:������b�Q޸�-2?�����ᆊ���]s�M�b�����IV�_ѫ9}G��P:6����C U�U|��t��/_�E�x�k�0���ub_{� 9K��)�S�"a,j�-9����]��4m�ړ6����[k��;�V�6[��<�������H���g�t������"�X�s,e�	#�a��=���YFL��Ф��!���з��� ;�t�,h[M��YZ�
4�������(�B)=�����9�4m��u�8���M'����h���q��eM$�����]>�}jI�K��c/p������� �(���������惟��� n�R� ���!;���S�-2j�����TYYm�!M7[�����r�g�VՕ�Om'���bO���������'���9
�"��F[���,�fO�JS�8x���?���v�U|�P�_@�~養���g2�O�'67���_�����^���y+1�Չ�w�Pz_��J�q�'
@5���z������I���,&|�"f��4���bX�hd~~ ��E�X�1����[?��K�g�"gϜ|��[�5{��J��	@�Z�� AMՆv$����� UI5F&m�����M����W�[_���N4"`w\�F|pb�d���U��弲��xWӿ�v�B�'&���B���~;Q�b���9kQ���4���g�����4	�?�[��Ć��M��M��'�"��oY��fc������^(���&�G��k��\���||U(��u�����]K��Q65�퍓^:� �DtZXY�ղ���xN"��q�+�ؽϨ�Y����=g���荥ٌ2�G�9r?Mys�x�kf�!�Ip���:~Vo��
���z?+���7�~� �@2��`�/~����Aܦ��y�n´�%$�]��H%��s�o�c��cz�t��b��������m4����!9��j��Z�H<���Q�90C⑐}n�X�D`�@ Z���	�,h��+5/�)��u��ib%h~�O~�����I�9�W����>�g`p���~���)���x��UOOO[��V�Po�y��$�I�R<���<��S�9��<��3���8�G�R#���
�eֳ�M3�B�H_�� ���� DXv)�­��M�Bj�J���� ��"�3@�V�����C�&����g�f2�AH��+y��W�34|�W_"O�0�F�Q�X,���o1��D$c|�O<��R���&���7�u�[$�2}�8�:�ًW(�J����,;�eE�[@{�",�4->��Pox�d��'�BWr+u�E�����߰���z�������~�k�p�g\�~?�9s�J&�$	 l���ٹ�o./-s��9j�*�T���z���~Ο��w��33s����{'�˝�6��!�U:�e�����X�V��>LՊ�hh�E�(�!���*��M̊��Z��?�O?�؞4Mg��8�X��gN���N��0�.]P�a��:*�������o����LLLp��Ì���^�/��/9y�$�02� �݋I��������5|!P��fE��b;���*�Ԣ0��>�����
������S���KN�z�W^~���sĢ+fs��!l��ݷ�fue���;�ҋ'q���Q̈M!_������~H�@?'N�����4�M<�ò,��2>>Αc�p��$3KY�W�7�D�I��aE����-{�S�3P�(�n��-"_)��XO?zҢ{t�WnL�ݿy�c&aItM�%������IΞ:&bȆ    IDATͥ˗�x�2�?�8�ϟ�N&�����o�ۜ9{�����O�ۿ�?G����O^�0�������aF�9}k��o�	�fQwX�P���}��)��¾f�k����G2�R*�ߕ�T.0;7˷��_��G���}�D����~���s{�7�_giq��O>��L��h�O���K��֛d��&�CCy�aNL�+fy�7x��u���>ҙ���,,,�Mץ�x��O_XH�A�"I�~%LI���=8���?�C�I$�ؑ�M�:��ɴ�#�������������`n%K��S$��8!�ҍP�YH�B9h�V$Z�-U
!�lc0���R;XQ��Δ��Z��~?����Ҩm:h)�̨P� ��G)|�k�|�d*N,E�ǏE�?{���
���O��4�4|��M��<�Z���66���r�J%&'��#��;��t:����/����3���24<J$�&�ƶ3�j>���4]E��"37BGI�5Z뙆�Y��B�	��[j`�:����7���z�D�Z!�͒�'�֫�?p��L7ÃCt�tS�ո}�.�K�LݺI>_`aq���5J�2�Z�ѽ���7�����Fc��'���}�ٻs8M������y��4����=��FݶQ�B�ua'3x@�RC�&��()	�B	�ZB
MJt-Խ(�R��#�-��G"a�+�Y���K�R�W��#��z���g��anܸ���9�7����Q,�y��7����A2�b��G�=��O<�aZ������g����k }=CD����{�@h��p�Ս_!��L7ʴ�5_��Jl���Y1l�
�|���
�O��'p"�I&��%ѨA�Z����\<�0��7�eGHg��tu�����kW�f�����Y[[eC4�}�9���0<����E���x�g/P�7B`E��G�S�-mpwaG��&�,�XM�h��M~%�1�MvװcL�+�-t�j� �K�T�ɇ�Ƣ�Y<�emu�t2�ѣ)V�4�&����;0�纬g7���'�Jp��%�\�L�X�Çy�'8z��d�����������q��9�׾��=Ź��9s�
�2�.��~.O
�����������5rs/j����
�#{�3����UT��ƕ�hJQ�T��Π ۶�d��;���/�����:�Z�L��'�~��O��ȑG I2jbh���y���A�m����>�=���\�5��F�X1�M�M������m?P�C���DZ�a�:��œO<J6�����15P��$���R.�A���0�������!�HQ�VYY]�\)S,Wq=��L7���_����m�w9�<��.�R����������k7XXY�O���g�_��$�C�6�CZ���s�Y��:�`KrhS'�� v���`���}��l]���{w��T�\� M���}4�%�{|��呇������������vJP;ֱP�X�vϾ����g�	�A�᱖�P�9���@hH�D3t�@)��b�L�H��t26#�bۑ{��PlC�uP�Pd����!�@� �o���\\��m[�Qbv��F�F�A����˯��^a��~��(��=�R��x�`hx��c{y��y��GH�2d2]��믿�7��_Pȗy≧XZɒ�b�I,;�n'Y[/Qs43��m�F�m|)QRC!��[�K�PB���@�4h��K)����1Mdye�����3�8Ϗ��'ܸ9�މ$�)�3]���clt/]]]D�===D"Q���رGx��SL�dbt�J���s����׮]���;���o��}�H${���W��[E7bX�$���R=hV���Ri6��Vc	�j�m��4�a�8�̮L�z���z!�Fl� ��,��2G�=ě��ɏ�3�]����9y�1��s`r���~�h�F���D8r��>��L�%�'���%~�������N�B'���׿��������wN1=�@�q�0���0c	\C��,���6�ȐB�1Z�eR�d��W�Bx>���lӦ�����eʥ{�G)�
�9w���EL3��:]��t���gl��²#�+U"f�����7�eGp=��+S<�����')���������0���2�f�)6|���M43���H���Xm}��'�����cԅ��98-�����������,'N� �N����:gϞ���M�ٳChR��d�T:����q��O��
�e��M)�Zo�/��s��y�8L�� =ü��)�9s��|�dw?�����􍎒-U�4_��Z�pó�ڹD{���+V�9����38La}CH^��IΞy��W��?<Hww/�a�hz���q��$J	_1y� �{��Ju��'�JR��q\��r����:�r��C�7����1*~���nq��V<�4c��q}�H4�P�Ž�gPDy����xA��Ib�ɓO<���,��
��Ģ6�c4M.��H.�g~a�X<I:Ӎ�(Bj�0<<F"�$����Ǟ�1��F����2k��x�-FFF"�����(�0�z�&�{�q��o�{/���/���4�@�ZA��Dy��$����-�����>��mR~@�yhn��p��?�S�=_���Gg�����iǫ�X�~��S#б���s���=�̭�u޸p�ksk�næ��hݶ4/�� ����妁R���
3!.ܩ%����D�:+���lH��s�a/2��� PHp��f�^�^��1[c�+�p��}��4+e�V��_�K���^/�?����k<��q��$}=]$�I��*�c{�,,-�D�{w�����<�܋,.,���|�����N�=��*V�EfW6�y{�xf���QGB,V�%®��h�R?�&
ښaRHT��o6PN�R �LW&Jw:�p_7��(����e�z��d�o�O=���w������cH��z
9b�����2i66rԚ�3�:s��>��b���	��`�=�F��w�p{�.�j�E�ba$��C�	�4�@|!	�fY��b00P��!p	�n��!L�S'bH�zRϣ�[�+n8<����B������?�>��O���S�H�&�H#��R���8{�gϜE�u���H��I�S�"iF�Lr��].]�b-Wd|��j���:p�%�JS��܅�(J���ׄ@��K���|�YE4j4V��}EDjLN�'fX��V)�H$|�Lx�B2�oG=��C�I%b��;^(����L���ܾ}��~�{ܸy������Hi ���Ş�Ire�ūwY.�Pv�x� ŦO`X����+�(��~n� h*@S�G�7J%�ؠKױ�C��ғ��,�β�r����S'���<�<r����8����x�G�XĎؤ�ҩ�TMj�d��癞��W_��͛tez8|�(�t�3�/s��5�J#�F�N��8F4ES������R�$�~�ۯؚCM��|��I[R˯ћI��c�7����י�q��^�j|�S'���'801A����X�������;.���D����¥Kܙ�ˍ�w���c�Xfpt?�<�4v<C��Y\�p{��#m|���� @�c���l���� ��po��0�1�%��8�g����/�z�MΜ~���;h���Х��y8�:�f���~�d�ސ	��b�(��a�&�i�N����ܾ}���Y���S�ױ,�H$��&�����3�����k�X�o}�o)�|#���Pveظ�ћm�"1�{I�>���3�r�w��g[8h;e�_HtDx~���Dk�V��ܳί�Ɵ���?�x4�د�uz;���T:����a�X���	|�A�"/��t�!5-���@y^�O �0���uOdD�Vf�^�������@34�ґ�A��h��xe�ᡚ�k���R	+��$��9J�?��˼��+D"�x�H4$&�Q�Tx���	E�P�Vup���u6�M���uw�s�/s��-�n ��Z���D� ��V�W8�\%w�"A��*h��t������/�5��K j(=F��Z��`e�++y^y������_�u��0�?@�T`��-�z{�>C�������K\�r���営^���q�%���sܞ����$��(V�Di��Y*橺��a�:��&"�W �B����@���5�!�kh�6�$l�tO?�ZE��5��S�����������g��'�z��:��l˲h6]�<�z?0"I4M��ɰgl͈�����ͭRs|R�=�--�?2��3��(A e;ۦ�4�%=��(eXhB�\_�X��44����;<�މ���XY�	�F�V!_,��2���
/��&��t�0��R�8�C�V�R�Rw\
�Eꎇ,�9th������Z�wN]���[4E\���!����O�W��Kˮ]�)Qx�Ro�m����t�J��8}�
�&'�76Lfp�@z��59}���]ahh�ё=����� 8{�{��9��o�p��E.\����"!0t�T*���У\�r�w�8�B��3�8|������-2���Ԭ�Em��Z����.T8�~ ���-չ15K��C9�4�T�kN��:˭�f�~B1_ n�Y����t�����Ϯ���H~#K�����r��MV�W�s� �L}ㇰi�d�B�c)�g9Wőq|��
��B�4|�i�6��7"��b���f�\�%�HӕN�N�i6�ԫ5N�4t��>�>4+��JX�����<��
�i�J�H&�(�����m<_ëy��e<ף��"�/"����J�
	%�,�f��Ǥ?����z��ʚ�#�z	���VA�RH�g�H�X�RJC�Hdt�c�ر��uwg�F"��mS��5�(K�*�e�}o�JC)�����P��d J��{B���L"a]�O_nU�nj@m���.�q������8nۈC��M� _�:�G�%�&�e�_sq�&n��m�<������D,�H"��[D$�F���
Y�gf�׫X�AĎ�i��h6]�#�0�o�RGi,,�Ss�++L�ΰ���K!-�6Itw�=��R�J E�*�@��PD�?Q�t�
��V�Zj��Ӓ�����P���H��1<܋��t���Ts��w��L������� �L��L��Y�.]b~~���^VW�q}�d����$�����Ynݝ��A�0t���H� #jk�!����;��[Y�6�Rp!#�����X�^�Q�#�h�|K�C���
�j�j��+L|-B$f�l69u��u$�U�!����+e�8}�C�D���te�Y+6��;���冏fF�Eb$�&�&��υ��03���#�0#,�@�M,]g��O3u���*~2�����2fD��+E���;��9d�Wi4jKy���O�X��"��a,-��n���!�����0C�Ì��O�����\�|�b���"O��?��C����
��%�am9��yw�r��(a�G�4�M|�Gj7�橹M�G��q&����3ܹ{���"7o�������*�D���Sljl�+H�q��5fgf�5}�F��������䡇��D�c\��������]���]k�}�;ֽ5YdG�(J�eY��ݲ��n;Ai�?� ��_$0$� ��F�iO�l�lJE��b�y��g�kȇ��νE�F˶���Bթ{�9{Xk��y��}�wy��or81�0ޟ��v�'�}����y��ۣ�����OMx��ZU��s?�t�ˈ�����3�K�]��c�8=2���3���M���[���M��W�z(�,����<v�,��>��s��9|�co\rk{�{�����IEUUɲ�.,m�O��Ǥ�ĦY����u�b�Ge9��2�k�L��3�S9�3.�§>�ɓ'�{�.���
W�\ax0�:KQ�LXYs��)�����:^w1��ZG��3��7n���M�����i:�U���t�s����Q�c��k"�?0���HJm!#�>
ïGI�Tx|�٧Y_Z�Dgc1@q1�G1!���:��A/�О^�af#r�T��[���)cx��>��8ِѤ���*F�~V.j 1xRE���b�[�Ik��s�:���3��t�q�^�b<� �Nv�~�GQ�������n:���"o��.Ã)��y�gY]�����y�m^����P��pZCV����l�=�-���!��Jvy�5K>}6�^B�����h6��)#k�v4K�>K'V���^��0�;`ei����s���؅s|��/��~���ɷ���p�����<�Ɖ����O����_~�e����8ϘY��N)&�䙧.�������d�r,�w��nO]1U^aq����O=���o���'��)�����iɉ�e6�^�l�{[,��`��agg��,k���RX�8���&"���5�,�,�s:�h4���;\�y�y,���/}��8������J�uk�Se�y���:�(�"�p��o���E��Ͼ�w��O`}�����&��|��gy���Y[_b{�!7n���������+r�,���d�h8��/s��y$�ܾ{�͍M�N�������O�����y�]z�eή�����~�O��"g/=�k���nb�#(:� ���� {[�E�E����ݻMy�>�����V�x�c/q�O1y뭷�������k���n��\�~���n����st;}^|�EΞ9��s��^}�{\��&�S�(��d��y�^|
+��l�)�b��	�S�U�6*v2vhS��t)tξ��Wn����Ǟ�ș��X=e�d4&�[������uv�ȋ�"S�,���qp0D��S'���e��%Fcn�~��)nm0�A��U�]����A�G�ɣsT�-A�k'��֘���K(DS�c%Ò����dn���ʍ�����������l���SL�p��C&�	�N���� `��t:4��x��;��s�6�ф���oc�0����Kg���"=g�?zG2�n���~�ؓ�"�:K�4eT>}��y���E��� ���?�qb����\�M�{Ξ9�͇�9xW��c^ي~�wAITy\��B��r���Ao�n��-���M��F ��z>T+s�Z�����Q�D%��ņct���C�����(KKfA��{n��af`mu�n�؟.=�y.lܻ���zͥK�x��gq����o��|����.����z��:��pʟ��
o��6Y'#����`zK}t�@�Y�GI0c�*��3#�#(�X���u�D0N��Ԅ ���#˸��9��乧�gC��p�P3aeS؟����<%9�gx�3�ܹǸu�."�`i�w��������S/tV��{�E9���s<~�i�O���ܾ݇� �O�s��~�e�(ƪ��X���M-���S9����C�X˅����9}���U:++� �%���}VV�����z�j�D�'�7X�ؠ��Ұ�?���c��̠��L����K��������_��}���讯#d�9�[,��+�2:��[zf�����o}�����os�`��>�<���q�����7���'>F��a��Fֳ�q���زd6�bg%��KO]"�v�u���=d<��pĝ�Λ�k.�;�0��[_��|�3O<��û�o0.��4�I�0W�ms�Q��T�
X�S����;��c��l�bl&���U�ߺ˙�u.>v��~��>�'.P�&�Ǉ�ل��Jd��/=�)K��%����//#y���]���-�>x��o��/ct���CV�l�ٟ�'�{�)�޺ύkW��`�{�TV����Ik�_-�}���eX�YCg�����?����;�:��R�`su��gY?k�{���5J)�ܺ��.��U.��prc���b3����q�>[�c+ɰ��xlq���V\Cu'у}��7��(�">���L������v���P�e��,�`j����.��bXz�|�*7>��s�������Nu1�0��p�R
�]ƈ�u0A)A�"#D+����N���9��'9w�q>�q���U��ё�U%)��3O���TL�F%��=��$�R���m��֚���>x���St5�z    IDAT�Q�b,�(.�b�H��J���7x��-�݌~�`l��sp�J���+�R��'@q����dm�<��9���+z�������8�����pY����Mf˫��g�`SN��i��Z����s�+�N�"��Jˉ����Y^^B���'Y�8����[w�u�{{{��<���{wos��K�G��K,o��;y�W�:��K-
���L��o�5�;��t��v2dbJ)2S��g�����.>�1N��ڐk���2��O���C�D���*�nܺÝ��N�L�S&e��N�|�E~��N1X����e���Lʒ<+�	�Y�
T�c8� ���|���A9ap�~2b��3�`������������ll.���<w�):K�L�Sz�>+�k}\V����_��]���`�htHYv�'t�}��>����S_�2���_�Թ���������l�=��hD񷜯"[�3���?�/���r��<�{�
w0�����ë������7oR9�O�!�3Ο=���*�6Ob���jg��'O�u
�?|����ai������.�)����XU0�X9y����\|�c����w�*{�c�����o�
p�dF�3n���7�������%�s���}c(�?*�z��+�<~���:��t4ׯ��z��`�3�0���ʕkNO�x�ţɌ�R��.>����W8��en=��Ɲ�XB�A�n�Ky�;�	��0
+*(���Ҕ��1�}��'�9w�4K�>��GkM7/������^�y��-G#��C���G�^!�%��8��T�A���Y#�TP.~��Q�ZE��#�x�����,�)���xL����Nk-&
$˫�����K lnn��t(�2�|jLi0��h]!*$#E��3��Q�>�����7�z��갼���J���H��f�&!F�Q���3PL�"�u"*^w�B�����>X�ز��'?�I���J��������O����^�Ko��z%��xH��GY��Q.>�T����FP��Vu�y�p��*ꑅ��e|�;W�\ԣ{��s�L�>&�I�K���x��u
:��̂�x��wrƓ1"����շ��փ{,-u�n��%gNmrok�W��Ji&�1�X�<����!�Ν�,/�cf�p8�+!��ɸ��s|��_�s?�E�y��u��<�pb譝|��p���Su��Yj�,:��|�CN�8[2�c�P�՛�h��<h�Ȳ�L�ey���i�my��U&�)w���;AiE��p��= ҥT����g>�W�Wy�cO���W�q�6�񈼷����(M�=D}�]5��+W�8/��\�� �� �P�"��4��>��l��qo7G��`����KK�z}VV������tR��r��m��P�!�+�0���`�?s�����|��.?����!o��C��qr}&��}t�B��;�w�x���
֖,��dR�d��uqY��g?ά����px�Ս{lnn�?,9y‫��`�)��S��WO&�x�`�0��?b�%E�G��gyy�n����i�|�n>�ǫ�����wPY�����[�*Zcc����:�����s��Uf��� _N�Z(︷u��[��9�^���Ҁ��u�Wz��[ ��i��jJ���!��[7�V�Q�9 Y���3����~�������Ǎ�wQ����C?`:vg�`}�~��tե��!Z�u��.KKK�M��}� Z_[���Ӭ��3�B��0��������C��)��C�W$�bu$�����_�,�*$v_���HU"Db@3J!2ɱޱ�w�w��:K�W�\���Lif����*���!8��ؠ�cV�𪋥@��C���w���55�_[_k]�����g&�v��W^���[��*�m$C| �6�)�����Sq���⩟�o��#�?"Y�w�p�%�	d��+>Tz����ے"��`���_�2O<6X/��������;�V�W N���4�t�=��J��!ݰLD4�Ǿ9��ޤ�����@2qM�fy��J��?�sO����i
��.�,b�з6��+K�3�0>U6�~x�.;[[���Y��
o��+,/w���pf�Jz�ef����[\�t����o��Ͻ���|�޻z�譮�$�Q�G��Z����p��d���1:ǖo��L	6*�?���>�� ��'6�~��;��� Q����͛7)��ԩSL������N���u~����g��w�������������.�n����T����ZV��x�(�9y��Z�����Z G�Cv�#�X���FS��ݼ���A��^��xx���d\�j�9�����:��3�Y���K_��l�=�_��w��o~�	K�U�=�C>X*<�o_��ڀO���^��tyX:qgJ���tLW��l��dY��ޘ��^cuu��R�r�t:�4cJ�N�C�/�+lV�[Z�.yf3��z��կ����ͷn�����W/��p���9|�ᕠ\S}�u��x4\�JģS�8�N��8w��p��p�9<���X2z�3s�;w�q��p��E!������8��,Z��6�f3˸�q��Y.=�4�?�$��2�������w_�r����Ne8�"+0�a����ڴ'��Z��|����@w��(�q�ab�~�D�$�
��xo����s�J��:�~��k�S�\-p�w��
ᾩH�M�0NkJ�z���`�p����������(�vvY]]Ɩe�˕�ݼW�F�^���|X>Я��\�q;����3�.�����
2�QY��x�A�TY���K�E���Ϛ�G���?�@�F�c5�*�:O9�Pt��t1%/}�i�,���X�����Q\���׮����/��mn�lq�i����,��^���`�G�4�%fm�R`
Z|0��Fy0F3�#$��W*V�����`����WV���b3T�ȜÔSTY�J�ì�`��J<��Z�!�
h��� Omn��p��dB�w޹�>g�|�O|�~�?�5�n=���m^���\����Q:��t)�'�u�.�àEt8	 3�������gK�l2����(cP|� ��z��8�,'�s�wL&�Y��=��S|�������x���?����w��{��(��O��W����n���&.H�{O��<�83g�h��%f6az0B�����s���Dg��!���Լ����R�iY2�}�|c������O��:O\~�����ߺ�7os����Ӧt�)>Ǧ�����{�8O�OrDޅ�����صs�<�t��0��1�����d�������y#�H!�ZȲ�������_�+������0������������-t���V2f>YE�� R�PP��$�!*�%^���f3�L�� R��1>�x3��E#d^Т��C�O�xJ�l�uu�W�4XZat8f����?�	>��ϲ���dZ����[������J��@M��C�
ב��ՠ�	�M������i�h\�{*>����	9��ۜ/�8��X֧�Z���~?�*���sM��pH\�ޔ�r�9!vZ�a��.(�ڲ�H�+�hP�չ��Pώ�����<��Tut�ʛ(�OiN�uН>��E�.�����g���$g���Zac?���{~p|���G�"�4%Nµ��=��`�)�3,i�x�7�k_�����k|��������b,�O�XT��x��c��/���&w��k�:F���0�e&%:��Вa"u3Xb���"�� O28����x�x�*�GG��z��zH��n�El�-h�EwoK�,�r�33������ʏY|������r`�I�*z<�O~����/�ٗ^be}��ѐ��\��W_�死LJ���� �4"Y~Do�c�?��Y]�	@Dk	������b$���FLיaf3�l2�΃ϰ�Hҍ���bi����/��O��O��
���)�C�v�o��6?x�}�?|���X9�����l�λd:��Y�N�f"@�P��8JkC��J�լ�C�l9���4Pm�>eZgAe�C�Th��Z+���$�ހ�;�'.���.7l�`xȟ��2ww�E��C)AT=/!K >��f�*��}p�S��-���K���+ ڡ�.�
E^��3���J�38�P*%T�X���~#��]�N�����o�6_��/�����������o����tɘ�-
��ŒB;�>*�)_�g��*`��#��}4q�nA��̴�Āq�2 ��y��J��*eHt�U�JϹ�����S<��E��>xp����y�~P�T
HTu%��@�wG(��,5�A���Us��$$S}�k�*�b?]C�X�;�8Ncd�f�L�R��QI&�KXN�씰�����Ra�0�����N�y�꾤D��*��ƾ�U\7��GE�]�^,
�`��<��c^�
�U-#���pI<*&��j�6���v����J��W7UL^�6(�v
v�~�`m��gWW��Sgy��H\��X ��X��ױ.����{?�3\�{�k�Pv�r�V��������2yo�hb�����h�+����{A��+W+��%��r¼x�
�%Z�j�����#&/��C>��M�Ru,%
%>��!�	Y���Sl���r
6b1ܸ|��_A&ˑ���2V����g?�s��$��en=�����x��ؾyV�譝��\:u�<h����	��V���5�:��j���O�I0�/(��u4*ϰ���h�S �)�PD�рR>��,�ɲ�Ҹy�����+3^��+��WŃ��ځ<���z�XR! �)H��RB2/��9�I�@&1��U���($S�=`R`fA�c0.d�CqE!y �Jb+���XZ�#�������w8����f���k7>ǞeK���=�[����z+��LۀJ�*�p>V�55Xr�4>�x�B�=�S�5���c���B �x���p�k�O������r탛|��pt�M��Eu
������ҤZ����/Ǆ֩B+�SF�6�c�(q����;���ҁu8Q(o�O��c�I'��Kws�ly��w������bo�.:HV �$z�����(}�׎v��W���ox<S���a��*P�C_�1��TW��ᪿ���׉��y�*dޯ��=魡QXD��`�ėJ�����������9?�\�؛=G�ٱ4e�
`��f���*ː���T�c��^���>�wAtH2c[W;��*YyD��#��޷���k\|���EP���������3��?�����S��sY��c1~B�bq/�?�q���g/���������`����ߧX������Oq8�L�%fj0�T�$U*R� �s�s��\�Yl ����h�ɰ�bM?OWA`��J;
OR�IA.Q��?�#��O�P�j���T��J����t�J 1~������f��'6x��1�q��-���)z]��k�.���NK����%��b�TPyIU);VE*�W���~��K*UP�P�J�CK�
� 䝵�fb�ޠT�"S
���(�3�B�����,��^xx�>�W��?s�\���y�`d[�,��I㾅ʴk$
�S&�
��)����W�+0�| �'�S�3Q
��X�M=t�yQ0�N�x�"w�����6�^�����ML�dJ�C�G�(B�#�:�F*���m�)>���fJ�I�Gpo�6�O�3����,C%
_<�J�NF��eyy�q���0�s�iɩ���R^I�WVA��G:��xU�\{�V��`?��&��Z�f�GE�o��PU��A�P��iqK`��H{��`um9��B���޽�����Y]�`2�8���oJ{W��\��<�	x{�.�}F�����֟4��1�鈽��u;�<��jn>�E��BDU4��c��
�C���N���h�&��0��U{`�f�ۊ�0��>��3w�EQ{^CB"E3V���� �:�r��X�PL�D[�<�{�1����#�\��E�G Ŵ?�9I�W�czgp�<v�<��p���\:���_�6�쟾D_x唖�.���X�P\���oܸ�������7���������`wj�J���&+�N�:}����݃��X����UWy��9�r�a��%�ן蝯�D4��M�����`���Ͱ>}����z�Ǯ�H��--88�dei���aƍEg�DtR��ͬA��-^2�4��A�k�
����D�m k�A_u��ub�+q�� �P�T1�N�9%B/�	��u[E��*�<�g����&�:�d>���zn�>$�w��hF/�M���h�Y%��|@q�җ^+U�)�+0�^I%��Rϓs��c��jW}kM00�gi��>�HN$� �s50sS���)$���f�c���s!�׊,R����јtx���+�}�i�	��@ݓ��?������c�GYOnHTQ�6�?���ޠ�\I�\J%$(������B%�e����b��XfN��8���5p�$��(��e"1YTq�u;�P�^EUS�@^��%�3p'�O2��s^w
YP��5������9���]��z.��w��W�~�B� Li��8K��.�O��[�\�5y,<L|�o��1�Y�G�GR3³$%�Tu׽sXo���J2;%wc�d����~�_��/q���3��v��b,�O�XPO��b|�s��-�������/ۻCT�!��ٔ��>32���A��(j�Rߦ�x��Ϛ=8ʵ�N݁K��C��み�j�h|�+)��Q���q��^e~<���&�Ƭ����� c,����nl�
 ȫ 4,>Rms��P���/����H���}╏Z�8K��J�%��OU[2TK��V&�� ?�u�}�8e.����:�_� �)�g(���g�Քa/A�K���
,k��ڏs�nL��U �@EG쒅�I1��&R�t����R�+�M�-"��UI�贠�^u���#t��*�m��(,��D�q[T�yOV���G�m��"�iv��tFGeXĉ̬�Ba<P/>�W�2k���D�L\?	��u�(|�mEޣ�&�y	@9���U-l�E���m���>�?!��]h�D�X��ڦ�+h���v$a��p
";����������l2�q�k���ժ��j�D�����{�����3	�MI�Ii�U¯�����D�� ^�W�/���\f]Q$��D(ĩ�.���佊t��+�)�e6��>
 ����`��Ϩ��J��x��iH�8�8�z����g>�)^x�iN�-S���p�z�,�b,��b,�?�x��������C��Ͼ͝�}lg�Ag��R�锱Ƈ:E��WP��iIa)i��;$����S@@������!f%IE��cA$�����u�w���^�Yϳ{�a��q�u^��5�rO	k��p]��(��F�E�rNj0�?HV�i�����2�L�q�B�b����8���>�t��>u�9M򞭪�aI�YU���o�>��9���I���#�
�c�T:ʢ帾�d�u��<��( Fs6Lo��n�����3�Tq���>�>Cl6��?%b��j�MgN.O9����e*o)��X�h��i�9<� ��)�d����
s�����
�����[L��_��K�b0�^F�q�I��kF�銏���V�g��zѢ�4e�<U�6:�AUՌZ��C��~�ncF��l]�6z���7�dᣴ�%g�9#����L�~�\�YzSn�\/S͂�B�Ő��R@y�E�^5aI�xٞ�m�)�9�M<v��{����'u�=��$����yН�������HY{����_G�#� �)O�@��m�(ITO`��8�-�9�@�tR�j`�v�f���wzY;I-����.>m��(�~�q��䄉�����>���v���G�>�G�p��?K{ѹ�7��!��ǰ����-����ep�K����H&��(���}����W��>t��mA��x���~�|���+PR-�VD��0���e�/���=����!v���ikM��r��
��/��0px��	į�qa��ȓT)I�1�"��l,ia�&��Ὕ尮�%�4">�Ҳ=�������E}��$�L�ͣ���G�~��, ��Xw6cˈƐ=K%�Ŭq7RH�4X�3P�0��d^S�9Ж|ɝ<����P5����HYm��|���R�%�f�Ɗ����[:�)�@�������I�˓?�埸������9�JZ�썋�}�=�|��_�G�C�21�b�y�P�s�/2�ܦo��_q�������q�����!��L)R�@Ml�(y��A9�o m�)r�����:{�-�t���:f�vb�и��F���0J��]��ys@�i*)�ӦU;�H[�@���by'k?�3�Km��	�������7�/BrU�TM�eM�6��-٨r�]�״���$��<m�Ւ2s6�=:��bW�Rק���Ǭ�[���1߶���yX�>�;,5�ʍX�s,�V7���@�ر>���|��ͺ&��e21��kG����{��y$�J�_?�-�mےvנz�<u���w��{,\�||�x��k��������]51��l��׼_=�a�O�u
w�T���>Zo~���b�VGg�2ac`K.x��������zEko>��f��i+&3K��8���T-1���]�?�;7W�|�`����%�fA)C�W�WK��H�(;���iT��g�ST�PxZ<��z���/+�zh�V�Zj�{J@�Q���=S�9jG�g�s=Ȩ�f������
-��U���=�ݱAM��J�;+}���H�)�n�!�.dp�h���c�M9Iy� ��oֿWm7�֨`�q�fJ:h�6]N�淓�x��b�"󟣷5��A/ܟ�3������h��<�;��h�F`"ޢ�?h=��3~���]��M�%�E#�,w�&��H��]��㬖f�a�H��-�GR �	1�d��$_�Q�7���W0��E���}�@�f�
X��N��(�JJ����-�N���r]0څ��0��8%�Z�V��}w��3�OJ��y������R��\w���{��0�+b��������:S�Լ�U�j�r-"��(X�m��6S�&)yߤo�a�N���T�.���Q���"��M�.^�Wc?
�e�d��;�I��V�N�8gP7���Q���[���?���pw�z}}/�U��9�'��o�R�2��d!0dx;'���1��UmGb����� �61��iN\^��&�"Ań9�^�a=9��U�%����(���b���Xm�;���*�Aŉ���n��5�x {��.k���Z������5s�ii_G�����cu�ז�O�}�-֨⺩G����D:`�/��<RV�iǗHEj5^#�_$�������s���v���	��t�����Sd��gs6R"��]\R"��`<�|��j��n��M����A^
%!��M�K-��17�kfߒ��X"C:n�"�Y
l�İi�A����d�*l���B�K�O��c:�M�rƃ�����hX=`��\{ �d��B?fo��w�T}ũ�f5�u�f�=���N����Z��3
]�6Ym�MνX��0ų8���,%����i��;��@NE��1֨�]��ߘ Z~Y!��|\�N?*ݑ8�ܘ�h��tHs>�&,e<
��=��A4zzO��B4��i�է�ݥ�@�"��鶫��]�N��w��Px�7Np�Ǝ��9I��1͟���N���fJ����G=e����r��L�8��ߜ�R�]$�4]�v	?��ѫ�9.�L���a/���]����F����/G��i۾9�L�w���L���,��~��o$�掱j2�;�"F#����;��7�%V��;�(�ɑ�Uԓ�D܋/�E+eh��K��1,\����g5x�FM[ϾJ
�5N��h���s)���=���ށ0�g�Ral�s��w�5r�7^� ��k��6Fݚ!�N��,�%��3~�]	P�J؉ˈmc`��^I�h��9�f�1����\^fSu_̀����R�WFVjr�\[�����l*.ۥ�� 2�	2�@�da�u��K�<��`�&�7E����b�bj���A���d m�J�c{�U�"�������uV�ee���n)�]QS��������.�]�����c<d������-�;�AnA���V�ܱ�k	ꉱ��B{?y�׈iZR���y�9+?�5��C���/#��ۦBTk�Z���,�M�W93�Hpm4���~�B��v����@��>�����߂��b��B��-�D����C#�E���C�'#��G����K���8d����ɑ�+�|Ľ�ixX�L�� c(d�u��vk��H���͍��^�}�hZ40edj��t>�\$�3���=��"�q����8�q�Ym�X�&�t7����,U��-����n�Oʵ�?�;�] ��`�y�"�H�0��O��I��x��������웊k����Wksʞ��]q��ly�zE��(�/V��Ե�RH���E?$A:����X�7�2�r"]lͪ�ŁV���Yҟ�({�������YC0�p�|W�qI��`QH�L*��a��
l_h�r�� 냳*�~F�*�$Ƃb��
��XC3B1Yc.:�o��:�����_�f���F�7Unf��Ɩ"KM����X�y���Z)l���OZ�Ro��63�A�[��Re,������
�Ɂ��m&�����Zʌ����0�pxG��nP �W���(��9�m����vz�R��C��[�8�%3�H�}r)yoW��5�i��b��r�r�E��ohDg��s)��
?o�S�O�Iw<.��B0(�EaF`�D��L������Nf,�N��(��OHd�e\����~k�����zf2!�-d��<�ɯް�B-���>���C�F�����򖷭�#�D�Iv�����}YHǦC��؈��Q��LZe�x�7���3j�9g�"�m��z��UO"��N�6�F�z8�Gw�[
�_[N,[�m�/)3�۝���y����/��	�?�4��CϮ{�o=��Z.�]ŏ�Y��f�A�B�m��1���0([ Դ��N��z�us懻�	���s����E�J���#�s �Ȕy�� jPXPh�f�������{�R���>"ct!X�(N"i~[�g�1��d���eKf��2ތE���eK<1@����E�?J����������"5�}��4m�(���->Z��Ġϵ����)���	��X]��c������������՚�b��J�ZB������QF�h��� ��{�2県�Zցuk��Ι{�H�Z��h�P_��������Ϙ�	$o꟯V�d�ض�cAL�/R��_63z�V]A?JZ�����JK��UP��zdxX2嘼�ݤ�ޝ9�m6Yy��N�΁���O���*�	d�����(Ҩ!���ho����	z����ɹJ�9K�ٰnz<��x��e��s�e��
�����S5\12��w7(ٽ��T(�)�#?�|r;v;ӹ�?s«�%�3��p�m����]WCO�8�Uǧ���p��[l]b���%�
�)ܘ��O[9:�.i�uf_ΌJ�|q���Cť�H�L����}��R)B&
đ!L�3Zk�k�L.�Cc=�b9;�͒�v�V�bW1��Q�D|lF��P$_`��{���fġ�ùgE�.�T�Y�"��$��1˄%\B�)�����2a�P�a_7�N����Fp͓O�;d�Ks�1G���Gb|�Fy 0��R�o`�*{dӥj�sJ���1��~��uqYiP�k��;�ųI*<�N�N��oG7�7i��v%�½�K�����@�ބT|����� yW�"�'�M���"ea ��79t}���ş8�R�����y��}o1E�E7<�{��[�c��멿���� :���x�Y�݃꒝���5�я��o�/�@��f�z��F�+�|�6[��R.��}>��1eaI��w�z�ԪL-��=������D����%���sq�g�#�~Һ���k�;��J��b6ʹ��bC�ѯ X�{ �,�=�;	[Er�tu~�i�-���w��t�2�����x=Dv#�q��94�Gz�B���T*�Dݜb{�xL�����ˡ��jVpݟ������������a�a��� ��]���,�p�_�>�Zj�Q����z����o��Q8�;��Oa�t�-�۠Z	OL������A<ts���BR} ��I�{�W��^'(a��F@�x�J#J_�g�0*˲��
L}g���c~ÌA,�_:O���ЦU�d�����3�Oq��T�CJ��߻ �L�.�~y�X���[�e�|�q����/t虄�7� �bn=��5�Ĝ����N�G*f<�`�� SV�،Z�I�>wC��-����&#�]�x�9�&�hɂ������_d(��-T��ro�mF�\a	Ֆ�$z��Ji��;��8��Z�Ty%��2�����=E� R݆��;ǩ��&D��X訕���G�z��/Ԃ��ݪ\rc8�Q��Ś���]��t�eJ$wi�E�#P/Uʌ��́�լ\��.����Rc�#�E�w3����v�Ը���6�MM�[��NZ���\Zcx��W��O�\ �?PJ�d��˿{\�vc��@��%�B��Ԅ.}��%�w�y�1�۲)!�����袹�����I�Ƶ���R������W�rS`�S��w�Ţ���0����� �ͪ&��%�I�B˕��xv{��d������a����\�����ꦎ��d��gK�4l�PS�#\kgw�'��H0�0�=v���ۨ����[�(��RV�� *�7af`�C�ZB�i*��3��R~�^]���3��P�>�d���Q\IT&�'G$�����?��$*���/��℡���_^E�F��)C9�;C9��WbC��*#*ă�a##�i���FN̹\��~Y�8�ǥm���9��:u�����ЕV�K�`8C�i��;��i@�^�"���N�)>	O[�yU6o��Hn&A�5��+�}�Е	�v0�=C]vb�p��+(���<\�"͎<ᓵMp
jԚ����58Mp(���B��)�A4r�v���j7 �i�O�FY��p�h�O�PM�����-�.����;�H��)�����zY��j��x;���O�Œ;�h�)���fsP�g,H��b��oK6jz����e�*��c���#�'B+�0j�g4�8ؠ��N����W�<�UC��K��8��~i��ѽ�7��7��$���}2���<�$
����|C`X���.��K�_q05�[���4�`���|��f��n�"��GV���G��U��)�o�k�z���x���o��F�_o�/HP���������8�9��ܛ�}�{vƩ�_��ҕ�ƫ��� Q�i��0�K�>�-�\)!���Iz<��K��2�L<��n��ɚAx�A�~M��&��ʌ�lx��m����9���a
�0�$ѳ;@��R��<_R�`T3$� rz$�L9����B��k� ��H�S�ߓȸ
�=��?�7l��I�(5�L5���ޔ+n�Rm"jI�Rl�#�\ޯq�t�<��Y��J�@&Z��t����6yZ&�S���l	��(��*��s�Y��f���f��%䋨6�O�k��u���_�C�8uN����,s�A���>L�������(LXg.����ws��Mԋ�a_^G*󉨞�+d�2���>9]�=>����F�"���J����y:��;&z}�iZ��z���v�^P��[q��_�Y���l�W����?v�L-�%�������=P�/'�D�u��q���,�٫�$�?%�O�)/��y�� ��6[F��1S�W�L�R��\J�w/���U��f���7��tn��RYKe��8{՚:E�&�&��<i���S����[8�`As*@�r�*��Kw8�����v��cn��0���q�-�˿��!/UKgP%ԡѧ7-�vv�V�g\�u:êcnbQ�4V���է����1}�ov�c_�T�1`%@@)��LB�����X�@�R�L�2B�����_c�0�g�vj�.����55�OT= �/IW�v�ĮC�Bylw�~�xnz<La�=�c�0{��a�������k]zk��r�&s��Q.%�Y�/�֊R�I�����'M���DXg?3<�9��o��l��2��H�+	M�S��a�|v�M鲪�4dXu�c2/Uq��*���ֵ-1�h�	�rY��ۉ0iff����~?x���|�/v<U�q��}�/����ӯ��͐jUWn��}�^kyJ�$_\u@Կ��������&o˿�H����D�+Y�'Ą��C����zP�i[����y�>`�"-QBiߒ>���m��d���_�)*�Q}�� Ȏ&�|dl���$� �����n�u�Ȝ�m��$gH�J9��D$}E��b�W$c�bmG�[ڕ����a�~~�̡��ܪ�1����Ε����Y.(V��S��������m��a��}����� ��!ȟ��*�D��1��w9�
ARkuzf��ci�aQIK �����:F�3��}(�8i��N�RDG�X��.J ds��q�hQs��n�Ke�_t���V���|�	�RZ��FO}���~-��m�A�K̬�X1�/�j��(i���@��v,n�b?fK�= C�b1v���RT�y�B��������D�SG{�K�A�Lq�fMV3��R��31뎻��}p�p��˾e���f�$G�ʅ���v���백:��	΍�l�m(��l�<f�!O�o��oi9�P�W��a�&�!�'Ny����nr<�5N:���p1Gb:XRA�"Z$�ӗ��S��B�o^�8��<��R�S�&�§i+� ���ץݒ�4�G�B���il�ܵ&�6b��X�[H�����b����* �h���Y6�B��1�!+5���+����Aӂ��n���h�&7X/�ڲ�F76���(ۇ6�MK��̭Bd�pU9�g�s��W�,>�QJeV�#ygQ�����G��%�=�1Zw��JV*�VӆO�vMn�2
�赅����n��[��r�x!��njN+�u�8v�@�=� OWly)g �C��Z�{�5��2�Q�&��n%�����C]7�b��Ɂq��Y�J�2<�7�v=����}�8o��˝~j4m��>�#��*�6���
��T�ËR���v��9�W���؞ncW[	�M���qޱz=�E_C�w�%��iP�r!��"ҟ���?be)���oN�t
��K?/|���p���W��ϻ#Nw�?5���{��m���3l�vVR.S��_Ɵ�-��������J��U
�Z�i����G�H5���~l�)�������,ʒ��'�B�G�?�M=R�l�W`��O գ%��_�X��>Iߣ�}�L�����0,{�����~��MVN���u���j�a�9�W�!�^��ů]�)&b��	p�:�>�(�?�y�
�5�6_	:ھQ��M�LW��:}��2��S__+�L��� �E�k?��zJ�mh>p����f$�O��+��#Ѯ-7�h�qLI���~����4-����5^h����h Y�L�{'��W����m�8�i����Q\���}�\��,H��=#0��wm��0���8:���E�4���;�-�ħKW��V�D�}��N�'0R���h<��Z��eW�Z�J�yܐ
�֦6���^��o4��t�TTj��G:�E;Y������h��&ǆ�����UY���S¼m�:��ybB�U�d�?�,���LNL�Vo#�fժHV�G�+��x��O{�/�G�<���|x���
<:qY튎ʛ9[��Qr��|���'���������}�7���wwy�w�Y��a��ִ�Ġ��5୏���Ea۠����/b����*�����������qT�d	���6�@t���a	J���+�̓-><���kU5����W�������yi�7W ��?c)l�Ns��� dMMo�c�O�!�6�j]5�;7Iy�Jn��-� �����GV�>����Sa=��Ʋó@S��WZn��s������4���(fO"
o/8�|������P�y�E�)�%�Gx���J]�6k���6{>W�F]P��+�dN&'����KB�c�}S��戏U=��������Vj��f���u��^Px�ܒ2f�P9��E��[��V63\�>��.��f~j�>n�uS��*�:��0+�R��Z=#�w�$I5H5&�]��9=��:j� YPf07��zH�.���&3l!x�A=����[�� y�����F'�bO����w�q��U�})�����Z��C��PK   c]WP(wi  6     jsons/user_defined.json��k�0���Y%�h�[i��acl�i�5�6q��+���^��o�������5ۚ����ג/��%r��F(	�c?��is;jP��;�ܳ���N�1B�'g~3wJa�mAW����ނ=�%������D	��A�C�%$<JY��a�z<J��q�X�Gi���X�rShQ7�ߓ�Q���k�]-�L.�vH��i��DU�3
b�bx`��{T�Co��� �/�J�ނ9+�-�sv@a�މ
*Q����!qGďN,C��,ޔ�qӊ��Σ��;�����%��9��Ʀ=v2;����q���������qޥ{#4�f%�j�qȱM`��9�������������PK   c]W����,  f�             ��    cirkitFile.jsonPK   c]W ��!�} $� /           ��Y  images/c261b03e-8211-44a8-b3b9-e5822ea41eae.pngPK   c]WP(wi  6             ���� jsons/user_defined.jsonPK      �   #�   